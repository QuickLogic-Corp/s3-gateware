/***************************************************
 Vendor        : QuickLogic Corp.
 File Name     : qlprim.v
 Description   : Behavioral model of Logic cell
 Revisions     : Added specify blocks for Logic cell, GPIO and RAM
 Author        : Kishor
*****************************************************/

// logic cell ------------------------------------------------------------------
`timescale 1ns/10ps
module P_LOGIC3 (
		 QST,
		 QDS,
		 TBS,
		 TAB,
		 TSL,
		 TA1,
		 TAS1,
		 TA2,
		 TAS2,
		 TB1,
		 TBS1,
		 TB2,
		 TBS2,
		 BAB,
		 BSL,
		 BA1,
		 BAS1,
		 BA2,
		 BAS2,
		 BB1,
		 BBS1,
		 BB2,
		 BBS2,
		 QDI,
		 QEN,
		 QCK,
		 QCKS,
		 QRT,
		 F1,
		 F2,
		 FS,
		 TZ,
		 CZ,
		 QZ,
		 FZ);
input QST;
input QDS;
input TBS;
input TAB;
input TA1;
input TAS1;
input TA2;
input TAS2;
input TB1;
input TBS1;
input TB2;
input TBS2;
input TSL;
input BAB;
input BSL;
input BA1;
input BAS1;
input BA2;
input BAS2;
input BB1;
input BBS1;
input BB2;
input BBS2;
input QDI;
input QEN;
input QCK;
input QCKS;
input QRT;
input F1;
input F2;
input FS;
output TZ;
output CZ;
output QZ;
output FZ;

wire TAI,TBI,BAI,BBI,TZI,BZI,CZI,QZI;
// wire declaration added by add_buf_port.pl (Tue Aug 30 15:15:38 2005)
wire QST_int ;
wire QDS_int ;
wire TBS_int ;
wire TAB_int ;
wire TA1_int ;
wire TAS1_int ;
wire TA2_int ;
wire TAS2_int ;
wire TB1_int ;
wire TBS1_int ;
wire TB2_int ;
wire TBS2_int ;
wire TSL_int ;
wire BAB_int ;
wire BSL_int ;
wire BA1_int ;
wire BAS1_int ;
wire BA2_int ;
wire BAS2_int ;
wire BB1_int ;
wire BBS1_int ;
wire BB2_int ;
wire BBS2_int ;
wire QDI_int ;
wire QEN_int ;
wire QCK_int ;
wire QCKS_int ;
wire QRT_int ;
wire F1_int ;
wire F2_int ;
wire FS_int ;
reg QZ_reg;


// buf instance for PORT delay added by add_buf_port.pl (Tue Aug 30 15:15:38 2005)
buf QST_buf (QST_int, QST) ;
buf QDS_buf (QDS_int, QDS) ;
buf TBS_buf (TBS_int, TBS) ;
buf TAB_buf (TAB_int, TAB) ;
buf TA1_buf (TA1_int, TA1) ;
buf TA2_buf (TA2_int, TA2) ;
buf TB1_buf (TB1_int, TB1) ;
buf TB2_buf (TB2_int, TB2) ;
buf TSL_buf (TSL_int, TSL) ;
buf BAB_buf (BAB_int, BAB) ;
buf BSL_buf (BSL_int, BSL) ;
buf BA1_buf (BA1_int, BA1) ;
buf BA2_buf (BA2_int, BA2) ;
buf BB1_buf (BB1_int, BB1) ;
buf BB2_buf (BB2_int, BB2) ;
buf QDI_buf (QDI_int, QDI) ;
buf QEN_buf (QEN_int, QEN) ;
buf QCK_buf (QCK_int, QCK) ;
buf QCKS_buf (QCKS_int, QCKS) ;
buf QRT_buf (QRT_int, QRT) ;
buf F1_buf (F1_int, F1) ;
buf F2_buf (F2_int, F2) ;
buf FS_buf (FS_int, FS) ;
buf TAS1_buf (TAS1_int, TAS1) ;
buf TAS2_buf (TAS2_int, TAS2) ;
buf TBS1_buf (TBS1_int, TBS1) ;
buf TBS2_buf (TBS2_int, TBS2) ;
buf BAS1_buf (BAS1_int, BAS1) ;
buf BAS2_buf (BAS2_int, BAS2) ;
buf BBS1_buf (BBS1_int, BBS1) ;
buf BBS2_buf (BBS2_int, BBS2) ;
initial
begin
	QZ_reg=1'b0;
end

assign TAP1 = TAS1_int ? ~TA1_int : TA1_int;  
assign TAP2 = TAS2_int ? ~TA2_int : TA2_int;
assign TBP1 = TBS1_int ? ~TB1_int : TB1_int;
assign TBP2 = TBS2_int ? ~TB2_int : TB2_int;
assign BAP1 = BAS1_int ? ~BA1_int : BA1_int; 
assign BAP2 = BAS2_int ? ~BA2_int : BA2_int; 
assign BBP1 = BBS1_int ? ~BB1_int : BB1_int; 
assign BBP2 = BBS2_int ? ~BB2_int : BB2_int; 
assign QCKP = QCKS_int ? QCK_int : ~QCK_int;

assign  TAI = TSL_int ? TAP2 : TAP1;   //changed here
assign  TBI = TSL_int ? TBP2 : TBP1;
assign  BAI = BSL_int ? BAP2 : BAP1;
assign  BBI = BSL_int ? BBP2 : BBP1;
assign  TZI = TAB_int ? TBI : TAI;
assign  BZI = BAB_int ? BBI : BAI;
assign  CZI = TBS_int ? BZI : TZI;
assign  QZI = QDS_int ? QDI_int : CZI;
assign  FZ = FS_int ? F2_int : F1_int;
assign TZ = TZI;
assign CZ = CZI;

assign QZ=QZ_reg;

/* synopsys translate off */
always @ (posedge QCKP)   
	if(~QRT_int && ~QST_int )
                if(QEN_int)
                  QZ_reg = QZI;
	
always @(QRT_int or QST_int)
	if(QRT_int)
		 QZ_reg = 1'b0;
	else if (QST_int)
		 QZ_reg = 1'b1;


/* synopsys translate_on */
/*********************************/

/***Logic Cell Specify Block Data***/

wire QEN_EQ_1_AN_QST_EQ_0_QCKS_0 = (QEN == 1'b1  && QST == 1'b0 && QCKS == 1'b0);
wire QEN_EQ_1_AN_QST_EQ_0_QCKS_1 = (QEN == 1'b1  && QST == 1'b0 && QCKS == 1'b1);
wire QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (QRT == 1'b0  && QST == 1'b0 && QCKS == 1'b0);
wire QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (QRT == 1'b0  && QST == 1'b0 && QCKS == 1'b1);
wire QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (QDS == 1'b1  && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (QDS == 1'b1  && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (QEN == 1'b1  && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (QEN == 1'b1  && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire QEN_EQ_1_AN_QRT_EQ_0_QCKS_0 = (QEN == 1'b1  && QRT == 1'b0 && QCKS == 1'b0);
wire QEN_EQ_1_AN_QRT_EQ_0_QCKS_1 = (QEN == 1'b1  && QRT == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b1  && BAB == 1'b1 && BSL == 1'b1 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b1  && BAB == 1'b1 && BSL == 1'b1 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b1  && BAB == 1'b1 && BSL == 1'b0 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b1  && BAB == 1'b1 && BSL == 1'b0 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b1  && BAB == 1'b0 && BSL == 1'b1 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b1  && BAB == 1'b0 && BSL == 1'b1 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b1  && BAB == 1'b0 && BSL == 1'b0 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b1  && BAB == 1'b0 && BSL == 1'b0 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b0  && TAB == 1'b1 && TSL == 1'b1 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b0  && TAB == 1'b1 && TSL == 1'b1 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b0  && TAB == 1'b1 && TSL == 1'b0 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b0  && TAB == 1'b1 && TSL == 1'b0 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b0  && TAB == 1'b0 && TSL == 1'b1 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b0  && TAB == 1'b0 && TSL == 1'b1 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b0  && TAB == 1'b0 && TSL == 1'b0 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b0  && TAB == 1'b0 && TSL == 1'b0 && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_0 = (TBS == 1'b0  && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_1 = (TBS == 1'b0  && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b0  && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b0  && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (TBS == 1'b1  && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (TBS == 1'b1  && QDS == 1'b0 && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
wire QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0 = (QDS == 1'b0  && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b0);
wire QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1 = (QDS == 1'b0  && QEN == 1'b1 && QRT == 1'b0 && QST == 1'b0 && QCKS == 1'b1);
specify

if ( TBS == 1'b1 && BAB == 1'b1 && BSL == 1'b1 && BBS2 == 1'b0 )
(BB2 => CZ) = (0,0);


if ( TBS == 1'b1 && BAB == 1'b1 && BSL == 1'b1 && BBS2 == 1'b1 )
(BB2 => CZ) = (0,0);


if ( TBS == 1'b1 && BAB == 1'b1 && BSL == 1'b0 && BBS1 == 1'b0 )
(BB1 => CZ) = (0,0);


if ( TBS == 1'b1 && BAB == 1'b1 && BSL == 1'b0 && BBS1 == 1'b1 )
(BB1 => CZ) = (0,0);


if ( TBS == 1'b1 && BAB == 1'b0 && BSL == 1'b1 && BAS2 == 1'b0 )
(BA2 => CZ) = (0,0);


if ( TBS == 1'b1 && BAB == 1'b0 && BSL == 1'b1 && BAS2 == 1'b1 )
(BA2 => CZ) = (0,0);


if ( TBS == 1'b1 && BAB == 1'b0 && BSL == 1'b0 && BAS1 == 1'b0 )
(BA1 => CZ) = (0,0);


if ( TBS == 1'b1 && BAB == 1'b0 && BSL == 1'b0 && BAS1 == 1'b1 )
(BA1 => CZ) = (0,0);


if ( TBS == 1'b0 && TAB == 1'b1 && TSL == 1'b1 && TBS2 == 1'b0 )
(TB2 => CZ) = (0,0);


if ( TBS == 1'b0 && TAB == 1'b1 && TSL == 1'b1 && TBS2 == 1'b1 )
(TB2 => CZ) = (0,0);


if ( TBS == 1'b0 && TAB == 1'b1 && TSL == 1'b0 && TBS1 == 1'b0 )
(TB1 => CZ) = (0,0);


if ( TBS == 1'b0 && TAB == 1'b1 && TSL == 1'b0 && TBS1 == 1'b1 )
(TB1 => CZ) = (0,0);


if ( TBS == 1'b0 && TAB == 1'b0 && TSL == 1'b1 && TAS2 == 1'b0 )
(TA2 => CZ) = (0,0);


if ( TBS == 1'b0 && TAB == 1'b0 && TSL == 1'b1 && TAS2 == 1'b1 )
(TA2 => CZ) = (0,0);


if ( TBS == 1'b0 && TAB == 1'b0 && TSL == 1'b0  && TAS1 == 1'b0 )
(TA1 => CZ) = (0,0);


if ( TBS == 1'b0 && TAB == 1'b0 && TSL == 1'b0 && TAS1 == 1'b1 )
(TA1 => CZ) = (0,0);


if ( TBS == 1'b0 )
(TSL => CZ) = (0,0);


if ( TBS == 1'b0 )
(TAB => CZ) = (0,0);


if ( TBS == 1'b1 )
(BSL => CZ) = (0,0);


if ( TBS == 1'b1 )
(BAB => CZ) = (0,0);


(TBS => CZ) = (0,0);

if ( TAB == 1'b1 && TSL == 1'b1 && TBS2 == 1'b0 )
(TB2 => TZ) = (0,0);


if ( TAB == 1'b1 && TSL == 1'b1 && TBS2 == 1'b1 )
(TB2 => TZ) = (0,0);


if ( TAB == 1'b1 && TSL == 1'b0 && TBS1 == 1'b0 )
(TB1 => TZ) = (0,0);


if ( TAB == 1'b1 && TSL == 1'b0 && TBS1 == 1'b1 )
(TB1 => TZ) = (0,0);


if ( TAB == 1'b0 && TSL == 1'b1 && TAS2 == 1'b0 )
(TA2 => TZ) = (0,0);


if ( TAB == 1'b0 && TSL == 1'b1 && TAS2 == 1'b1 )
(TA2 => TZ) = (0,0);


if ( TAB == 1'b0 && TSL == 1'b0 && TAS1 == 1'b0 )
(TA1 => TZ) = (0,0);


if ( TAB == 1'b0 && TSL == 1'b0 && TAS1 == 1'b1 )
(TA1 => TZ) = (0,0);


(TSL => TZ) = (0,0);

(TAB => TZ) = (0,0);

if ( FS == 1'b1 )
(F2 => FZ) = (0,0);


if ( FS == 1'b0 )
(F1 => FZ) = (0,0);


(FS => FZ) = (0,0);

(QRT => QZ) = (0,0);

(QCK => QZ) = (0,0);

if ( QCKS == 1'b1 )
(QCK => QZ) = (0,0);


(QST => QZ) = (0,0);

$removal (posedge QRT,posedge QST, 0);
$removal (negedge QRT,posedge QST, 0);


$recovery (posedge QRT,posedge QST, 0);
$recovery (negedge QRT,posedge QST, 0);


$removal( posedge QRT, negedge QCK &&& QEN_EQ_1_AN_QST_EQ_0_QCKS_0, 0);
$removal( negedge QRT, negedge QCK &&& QEN_EQ_1_AN_QST_EQ_0_QCKS_0, 0);


$removal( posedge QRT, posedge QCK &&& QEN_EQ_1_AN_QST_EQ_0_QCKS_1, 0);
$removal( negedge QRT, posedge QCK &&& QEN_EQ_1_AN_QST_EQ_0_QCKS_1, 0);


$recovery( posedge QRT, negedge QCK &&& QEN_EQ_1_AN_QST_EQ_0_QCKS_0, 0);
$recovery( negedge QRT, negedge QCK &&& QEN_EQ_1_AN_QST_EQ_0_QCKS_0, 0);


$recovery( posedge QRT, posedge QCK &&& QEN_EQ_1_AN_QST_EQ_0_QCKS_1, 0);
$recovery( negedge QRT, posedge QCK &&& QEN_EQ_1_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge QEN, negedge QCK &&& QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge QEN, negedge QCK &&& QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge QEN &&& QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge QEN &&& QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge QEN, posedge QCK &&& QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge QEN, posedge QCK &&& QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge QEN &&& QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge QEN &&& QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge QDI, negedge QCK &&& QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge QDI, negedge QCK &&& QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge QDI &&& QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge QDI &&& QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge QDI, posedge QCK &&& QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge QDI, posedge QCK &&& QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge QDI &&& QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge QDI &&& QDS_EQ_1_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge QDS, negedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge QDS, negedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge QDS &&& QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge QDS &&& QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge QDS, posedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge QDS, posedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge QDS &&& QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge QDS &&& QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$recovery( posedge QST, negedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_QCKS_0, 0);
$recovery( negedge QST, negedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_QCKS_0, 0);


$recovery( posedge QST, posedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_QCKS_1, 0);
$recovery( negedge QST, posedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_QCKS_1, 0);


$removal( posedge QST, negedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_QCKS_0, 0);
$removal( negedge QST, negedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_QCKS_0, 0);


$removal( posedge QST, posedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_QCKS_1, 0);
$removal( negedge QST, posedge QCK &&& QEN_EQ_1_AN_QRT_EQ_0_QCKS_1, 0);


$setup( posedge BB2, negedge QCK &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge BB2, negedge QCK &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge BB2 &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge BB2 &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge BB2, posedge QCK &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge BB2, posedge QCK &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge BB2 &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge BB2 &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge BB1, negedge QCK &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge BB1, negedge QCK &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge BB1 &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge BB1 &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge BB1, posedge QCK &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge BB1, posedge QCK &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge BB1 &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge BB1 &&& TBS_EQ_1_AN_BAB_EQ_1_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge BA2, negedge QCK &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge BA2, negedge QCK &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge BA2 &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge BA2 &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge BA2, posedge QCK &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge BA2, posedge QCK &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge BA2 &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge BA2 &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge BA1, negedge QCK &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge BA1, negedge QCK &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge BA1 &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge BA1 &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge BA1, posedge QCK &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge BA1, posedge QCK &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge BA1 &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge BA1 &&& TBS_EQ_1_AN_BAB_EQ_0_AN_BSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge TB2, negedge QCK &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge TB2, negedge QCK &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge TB2 &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge TB2 &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge TB2, posedge QCK &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge TB2, posedge QCK &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge TB2 &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge TB2 &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge TB1, negedge QCK &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge TB1, negedge QCK &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge TB1 &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge TB1 &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge TB1, posedge QCK &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge TB1, posedge QCK &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge TB1 &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge TB1 &&& TBS_EQ_0_AN_TAB_EQ_1_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge TA2, negedge QCK &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge TA2, negedge QCK &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge TA2 &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge TA2 &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge TA2, posedge QCK &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge TA2, posedge QCK &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge TA2 &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge TA2 &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge TA1, negedge QCK &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge TA1, negedge QCK &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge TA1 &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge TA1 &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge TA1, posedge QCK &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge TA1, posedge QCK &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge TA1 &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge TA1 &&& TBS_EQ_0_AN_TAB_EQ_0_AN_TSL_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge TSL, negedge QCK &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_0, 0);
$setup( negedge TSL, negedge QCK &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_0, 0);


$hold( negedge QCK, posedge TSL &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_0, 0);
$hold( negedge QCK, negedge TSL &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_0, 0);


$setup( posedge TSL, posedge QCK &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_1, 0);
$setup( negedge TSL, posedge QCK &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_1, 0);


$hold( posedge QCK, posedge TSL &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_1, 0);
$hold( posedge QCK, negedge TSL &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_EQ_1, 0);


$setup( posedge TAB, negedge QCK &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge TAB, negedge QCK &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge TAB &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge TAB &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge TAB, posedge QCK &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge TAB, posedge QCK &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge TAB &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge TAB &&& TBS_EQ_0_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge BSL, negedge QCK &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge BSL, negedge QCK &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge BSL &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge BSL &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge BSL, posedge QCK &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge BSL, posedge QCK &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge BSL &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge BSL &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge BAB, negedge QCK &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge BAB, negedge QCK &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge BAB &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge BAB &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge BAB, posedge QCK &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge BAB, posedge QCK &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge BAB &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge BAB &&& TBS_EQ_1_AN_QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$setup( posedge TBS, negedge QCK &&& QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$setup( negedge TBS, negedge QCK &&& QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$hold( negedge QCK, posedge TBS &&& QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);
$hold( negedge QCK, negedge TBS &&& QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_0, 0);


$setup( posedge TBS, posedge QCK &&& QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$setup( negedge TBS, posedge QCK &&& QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


$hold( posedge QCK, posedge TBS &&& QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);
$hold( posedge QCK, negedge TBS &&& QDS_EQ_0_AN_QEN_EQ_1_AN_QRT_EQ_0_AN_QST_EQ_0_QCKS_1, 0);


endspecify

/***********************************/

/***********************************/
endmodule    


`timescale 1ns/10ps

module P_BIDIR3 (	
		ESEL,
		IE,
		OSEL,
		OQI,
		OQE,	
		DS,
		FIXHOLD,
		IZ,
		IQZ,
		IQE,
		IQC,
		IQCS,
		IQR,
		WPD,
		INEN,
		IQIN,
		IP
		);
				
input ESEL;
input IE;
input OSEL;
input OQI;
input OQE;
input DS;
input FIXHOLD;
output IZ;
output IQZ;
input IQE;
input IQC;
input IQCS;
input INEN;
input IQIN;
input IQR;
input WPD;
inout IP;

reg EN_reg, OQ_reg, IQZ;
wire rstn, EN, OQ, AND_OUT, IQCP;

wire FIXHOLD_int;	
wire ESEL_int;
wire IE_int;
wire OSEL_int;
wire OQI_int;
wire DS_int;
wire INEN_int;
wire OQE_int;
wire IQE_int;
wire IQC_int;
wire IQCS_int;
wire IQR_int;
wire WPD_int;

parameter IOwithOUTDriver = 0;        //  has to be set for IO with out Driver

buf IQIN_buf (IQIN_int,IQIN);	
buf FIXHOLD_buf (FIXHOLD_int,FIXHOLD);	
buf WPD_buf (WPD_int,WPD);
buf DS_buf (DS_int,DS);
buf INEN_buf (INEN_int,INEN);
buf IQC_buf (IQC_int,IQC);
buf IQCS_buf (IQCS_int,IQCS);
buf IQR_buf (IQR_int,IQR);
buf ESEL_buf (ESEL_int,ESEL);
buf IE_buf (IE_int,IE);
buf OSEL_buf (OSEL_int,OSEL);
buf OQI_buf (OQI_int,OQI);
buf OQE_buf (OQE_int,OQE);
buf IQE_buf (IQE_int,IQE);

assign rstn = ~IQR_int;
assign IQCP = IQCS_int ? ~IQC_int : IQC_int;
 if (IOwithOUTDriver)
 begin
	assign AND_OUT = IQIN_int;

	assign IZ = IP;
 end
 else
  begin
	assign AND_OUT = INEN_int ? IP : 1'b0;

	assign IZ = AND_OUT;
 end
assign EN = ESEL_int ? IE_int : EN_reg ;

assign OQ = OSEL_int ? OQI_int : OQ_reg ;

assign IP = EN ? OQ : 1'bz;

assign (highz1,pull0) IP = WPD ? 1'b0 : 1'b1;
initial
	begin		
		//Power on reset
		EN_reg	= 1'b0;
		OQ_reg= 1'b0;
		IQZ=1'b0;
	end
always @(posedge IQCP or negedge rstn)
	if (~rstn)
		EN_reg <= 1'b0;
	else
		EN_reg <= IE_int;

always @(posedge IQCP or negedge rstn)
	if (~rstn)
		OQ_reg <= 1'b0;
	else
		if (OQE_int)
			OQ_reg <= OQI_int;
			
			
always @(posedge IQCP or negedge rstn)		
	if (~rstn)
		IQZ <= 1'b0;
	else
		if (IQE_int)
			IQZ <= AND_OUT;
		
wire gpio_c18 = (OSEL == 1'b1  && IE == 1'b1 && IQE == 1'b1 && FIXHOLD == 1'b1 && DS == 1'b1 && IQCS == 1'b1);
wire gpio_c16 = (OSEL == 1'b1  && IE == 1'b1 && IQE == 1'b1 && FIXHOLD == 1'b1 && DS == 1'b0 && IQCS == 1'b1);
wire gpio_c14 = (OSEL == 1'b1  && IE == 1'b1 && IQE == 1'b1 && FIXHOLD == 1'b0 && DS == 1'b1 && IQCS == 1'b1);
wire gpio_c12 = (OSEL == 1'b1  && IE == 1'b1 && IQE == 1'b1 && FIXHOLD == 1'b0 && DS == 1'b0 && IQCS == 1'b1);
wire gpio_c10 = (OSEL == 1'b0  && OQE == 1'b1 && IQCS == 1'b1);
wire gpio_c8 = (OSEL == 1'b1  && IE == 1'b1 && IQE == 1'b1 && FIXHOLD == 1'b1 && DS == 1'b1 && IQCS == 1'b0);
wire gpio_c6 = (OSEL == 1'b1  && IE == 1'b1 && IQE == 1'b1 && FIXHOLD == 1'b1 && DS == 1'b0 && IQCS == 1'b0);
wire gpio_c4 = (OSEL == 1'b1  && IE == 1'b1 && IQE == 1'b1 && FIXHOLD == 1'b0 && DS == 1'b1 && IQCS == 1'b0);
wire gpio_c2 = (OSEL == 1'b1  && IE == 1'b1 && IQE == 1'b1 && FIXHOLD == 1'b0 && DS == 1'b0 && IQCS == 1'b0);
wire gpio_c0 = (OSEL == 1'b0  && OQE == 1'b1 && IQCS == 1'b0);
wire gpio_c30 = (IQE == 1'b1  && FIXHOLD == 1'b1 && INEN == 1'b1 && IQCS == 1'b1);
wire gpio_c28 = (IQE == 1'b1  && FIXHOLD == 1'b0 && INEN == 1'b1 && IQCS == 1'b1);
wire gpio_c22 = (IQE == 1'b1  && FIXHOLD == 1'b1 && INEN == 1'b1 && IQCS == 1'b0);
wire gpio_c20 = (IQE == 1'b1  && FIXHOLD == 1'b0 && INEN == 1'b1 && IQCS == 1'b0);
specify
if ( IQE == 1'b1  )
(IQC => IQZ) = (0,0,0,0,0,0);
(IQR => IQZ) = (0,0);
if ( IE == 1'b1 && OQE == 1'b1  )
(IQC => IZ) = (0,0,0,0,0,0);
//if ( IE == 1'b0 )
//(IP => IZ) = (0,0);
if ( IE == 1'b0 && INEN == 1'b1  )
(IP => IZ) = (0,0);
$setup (posedge IE,negedge IQC, 0);
$setup (negedge IE,negedge IQC, 0);
$hold (negedge IQC,posedge IE, 0);
$hold (negedge IQC,negedge IE, 0);
$setup (posedge IE,posedge IQC, 0);
$setup (negedge IE,posedge IQC, 0);
$hold (posedge IQC,posedge IE, 0);
$hold (posedge IQC,negedge IE, 0);
$setup( posedge OQI, negedge IQC &&& gpio_c18, 0);
$setup( negedge OQI, negedge IQC &&& gpio_c18, 0);
$hold( negedge IQC, posedge OQI &&& gpio_c18, 0);
$hold( negedge IQC, negedge OQI &&& gpio_c18, 0);
$setup( posedge OQI, negedge IQC &&& gpio_c16, 0);
$setup( negedge OQI, negedge IQC &&& gpio_c16, 0);
$hold( negedge IQC, posedge OQI &&& gpio_c16, 0);
$hold( negedge IQC, negedge OQI &&& gpio_c16, 0);
$setup( posedge OQI, negedge IQC &&& gpio_c14, 0);
$setup( negedge OQI, negedge IQC &&& gpio_c14, 0);
$hold( negedge IQC, posedge OQI &&& gpio_c14, 0);
$hold( negedge IQC, negedge OQI &&& gpio_c14, 0);
$setup( posedge OQI, negedge IQC &&& gpio_c12, 0);
$setup( negedge OQI, negedge IQC &&& gpio_c12, 0);
$hold( negedge IQC, posedge OQI &&& gpio_c12, 0);
$hold( negedge IQC, negedge OQI &&& gpio_c12, 0);
$setup( posedge OQI, negedge IQC &&& gpio_c10, 0);
$setup( negedge OQI, negedge IQC &&& gpio_c10, 0);
$hold( negedge IQC, posedge OQI &&& gpio_c10, 0);
$hold( negedge IQC, negedge OQI &&& gpio_c10, 0);
$setup( posedge OQI, posedge IQC &&& gpio_c8, 0);
$setup( negedge OQI, posedge IQC &&& gpio_c8, 0);
$hold( posedge IQC, posedge OQI &&& gpio_c8, 0);
$hold( posedge IQC, negedge OQI &&& gpio_c8, 0);
$setup( posedge OQI, posedge IQC &&& gpio_c6, 0);
$setup( negedge OQI, posedge IQC &&& gpio_c6, 0);
$hold( posedge IQC, posedge OQI &&& gpio_c6, 0);
$hold( posedge IQC, negedge OQI &&& gpio_c6, 0);
$setup( posedge OQI, posedge IQC &&& gpio_c4, 0);
$setup( negedge OQI, posedge IQC &&& gpio_c4, 0);
$hold( posedge IQC, posedge OQI &&& gpio_c4, 0);
$hold( posedge IQC, negedge OQI &&& gpio_c4, 0);
$setup( posedge OQI, posedge IQC &&& gpio_c2, 0);
$setup( negedge OQI, posedge IQC &&& gpio_c2, 0);
$hold( posedge IQC, posedge OQI &&& gpio_c2, 0);
$hold( posedge IQC, negedge OQI &&& gpio_c2, 0);
$setup( posedge OQI, posedge IQC &&& gpio_c0, 0);
$setup( negedge OQI, posedge IQC &&& gpio_c0, 0);
$hold( posedge IQC, posedge OQI &&& gpio_c0, 0);
$hold( posedge IQC, negedge OQI &&& gpio_c0, 0);
$setup (posedge OQE,negedge IQC, 0);
$setup (negedge OQE,negedge IQC, 0);
$hold (negedge IQC,posedge OQE, 0);
$hold (negedge IQC,negedge OQE, 0);
$setup (posedge OQE,posedge IQC, 0);
$setup (negedge OQE,posedge IQC, 0);
$hold (posedge IQC,posedge OQE, 0);
$hold (posedge IQC,negedge OQE, 0);
$setup (posedge IQIN,negedge IQC, 0);
$setup (negedge IQIN,negedge IQC, 0);
$hold (negedge IQC,posedge IQIN, 0);
$hold (negedge IQC,negedge IQIN, 0);
$setup (posedge IQIN,posedge IQC, 0);
$setup (negedge IQIN,posedge IQC, 0);
$hold (posedge IQC,posedge IQIN, 0);
$hold (posedge IQC,negedge IQIN, 0);
$setup (posedge IQE,negedge IQC, 0);
$setup (negedge IQE,negedge IQC, 0);
$hold (negedge IQC,posedge IQE, 0);
$hold (negedge IQC,negedge IQE, 0);
$setup (posedge IQE,posedge IQC, 0);
$setup (negedge IQE,posedge IQC, 0);
$hold (posedge IQC,posedge IQE, 0);
$hold (posedge IQC,negedge IQE, 0);
$recovery (posedge IQR,negedge IQC, 0);
$recovery (negedge IQR,negedge IQC, 0);
$removal (posedge IQR,negedge IQC, 0);
$removal (negedge IQR,negedge IQC, 0);
$recovery (posedge IQR,posedge IQC, 0);
$recovery (negedge IQR,posedge IQC, 0);
$removal (posedge IQR,posedge IQC, 0);
$removal (negedge IQR,posedge IQC, 0);
$setup( posedge IP, negedge IQC &&& gpio_c30, 0);
$setup( negedge IP, negedge IQC &&& gpio_c30, 0);
$hold( negedge IQC, posedge IP &&& gpio_c30, 0);
$hold( negedge IQC, negedge IP &&& gpio_c30, 0);
$setup( posedge IP, negedge IQC &&& gpio_c28, 0);
$setup( negedge IP, negedge IQC &&& gpio_c28, 0);
$hold( negedge IQC, posedge IP &&& gpio_c28, 0);
$hold( negedge IQC, negedge IP &&& gpio_c28, 0);
$setup( posedge IP, posedge IQC &&& gpio_c22, 0);
$setup( negedge IP, posedge IQC &&& gpio_c22, 0);
$hold( posedge IQC, posedge IP &&& gpio_c22, 0);
$hold( posedge IQC, negedge IP &&& gpio_c22, 0);
$setup( posedge IP, posedge IQC &&& gpio_c20, 0);
$setup( negedge IP, posedge IQC &&& gpio_c20, 0);
$hold( posedge IQC, posedge IP &&& gpio_c20, 0);
$hold( posedge IQC, negedge IP &&& gpio_c20, 0);
(IE => IP) = (0,0,0,0,0,0);
if ( IE == 1'b1 )
(OQI => IP) = (0,0);
(IQC => IP) = (0,0,0,0,0,0);
if ( IE == 1'b1 && OQE == 1'b1  )
(IQC => IP) = (0,0,0,0,0,0);
if ( IE == 1'b0 )
(IQR => IP) = (0,0);
endspecify
endmodule

//-------- RAM -----------

`timescale 1ns/10ps
//pragma synthesis_off
module fifo_controller_model(
	 Rst_n,
	 Push_Clk,
	 Pop_Clk,
	
	 Fifo_Push,
	 Fifo_Push_Flush,
	 Fifo_Full,
	 Fifo_Full_Usr,
	
	 Fifo_Pop,
	 Fifo_Pop_Flush,
	 Fifo_Empty,
	 Fifo_Empty_Usr,
	
	 Write_Addr,
	
	 Read_Addr,
	 												 
	 //	 Static Control Signals
	 Fifo_Ram_Mode,
	 Fifo_Sync_Mode,
	 Fifo_Push_Width,
	 Fifo_Pop_Width
	  );

	

  //************* PPII 4K Parameters **************************//
	
  parameter MAX_PTR_WIDTH   = 12;
  
  parameter DEPTH1 = (1<<(MAX_PTR_WIDTH-3));
  parameter DEPTH2 = (1<<(MAX_PTR_WIDTH-2));
  parameter DEPTH3 = (1<<(MAX_PTR_WIDTH-1));
  
  parameter D1_QTR_A = MAX_PTR_WIDTH - 5;
  parameter D2_QTR_A = MAX_PTR_WIDTH - 4;
  parameter D3_QTR_A = MAX_PTR_WIDTH - 3;

	
	input	Rst_n;
	input	Push_Clk;
	input	Pop_Clk;
	
	input	Fifo_Push;
	input	Fifo_Push_Flush;
	output	Fifo_Full;
	output	[3:0]  Fifo_Full_Usr;
                            		
	input	Fifo_Pop;
	input	Fifo_Pop_Flush;
	output	Fifo_Empty;
	output	[3:0]  Fifo_Empty_Usr;
	
	output	[MAX_PTR_WIDTH-2:0]  Write_Addr;
	
	output	[MAX_PTR_WIDTH-2:0]  Read_Addr;
		
	input  Fifo_Ram_Mode;
	input  Fifo_Sync_Mode;
	input  [1:0] Fifo_Push_Width;
	input  [1:0] Fifo_Pop_Width;
	
	reg    flush_pop_clk_tf;
	reg    flush_pop2push_clk1;
	reg    flush_push_clk_tf;
	reg    flush_push2pop_clk1;
	reg    pop_local_flush_mask;
	reg    push_flush_tf_pop_clk;
	reg    pop2push_ack1;
	reg    pop2push_ack2;
	reg    push_local_flush_mask;
	reg    pop_flush_tf_push_clk;
	reg    push2pop_ack1;
	reg    push2pop_ack2;
	
	reg    fifo_full_flag_f;
	reg    [3:0]  Fifo_Full_Usr;

	reg    fifo_empty_flag_f;
	reg    [3:0]  Fifo_Empty_Usr;

	reg    [MAX_PTR_WIDTH-1:0]  push_ptr_push_clk;
	reg    [MAX_PTR_WIDTH-1:0]  pop_ptr_push_clk;
	reg    [MAX_PTR_WIDTH-1:0]  pop_ptr_async;	    
	reg    [MAX_PTR_WIDTH-1:0]  pop_ptr_pop_clk ;
	reg    [MAX_PTR_WIDTH-1:0]  push_ptr_pop_clk;
	reg    [MAX_PTR_WIDTH-1:0]  push_ptr_async;

	reg    [1:0]  push_ptr_push_clk_mask;
	reg    [1:0]  pop_ptr_pop_clk_mask;

	reg    [MAX_PTR_WIDTH-1:0]  pop_ptr_push_clk_mux;
	reg    [MAX_PTR_WIDTH-1:0]  push_ptr_pop_clk_mux;

	reg    match_room4none;		
	reg    match_room4one;		
	reg    match_room4half;  	      
	reg    match_room4quart;

	reg    match_all_left;
	reg    match_half_left;
	reg    match_quart_left;

 	reg   [MAX_PTR_WIDTH-1:0]   depth1_reg;
 	reg   [MAX_PTR_WIDTH-1:0]   depth2_reg;
 	reg   [MAX_PTR_WIDTH-1:0]   depth3_reg;
  

	wire	push_clk_rst;
	wire	push_clk_rst_mux;
	wire	push_flush_done;
	wire	pop_clk_rst;
	wire	pop_clk_rst_mux;
	wire	pop_flush_done;

	wire	push_flush_gated;
	wire	pop_flush_gated;
	                          	
	wire	[MAX_PTR_WIDTH-2:0] Write_Addr;
	wire	[MAX_PTR_WIDTH-2:0] Read_Addr;
	
	wire	[MAX_PTR_WIDTH-1:0] push_ptr_push_clk_plus1;
	wire	[MAX_PTR_WIDTH-1:0] next_push_ptr_push_clk;
	wire	[MAX_PTR_WIDTH-1:0] pop_ptr_pop_clk_plus1;
	wire	[MAX_PTR_WIDTH-1:0] next_pop_ptr_pop_clk;
	wire	[MAX_PTR_WIDTH-1:0] next_push_ptr_push_clk_mask;
	wire	[MAX_PTR_WIDTH-1:0] next_pop_ptr_pop_clk_mask;

	wire	[MAX_PTR_WIDTH-1:0] pop_ptr_push_clk_l_shift1;
	wire	[MAX_PTR_WIDTH-1:0] pop_ptr_push_clk_l_shift2;
	wire	[MAX_PTR_WIDTH-1:0] pop_ptr_push_clk_r_shift1;
	wire	[MAX_PTR_WIDTH-1:0] pop_ptr_push_clk_r_shift2;

	wire	[MAX_PTR_WIDTH-1:0] push_ptr_pop_clk_l_shift1;
	wire	[MAX_PTR_WIDTH-1:0] push_ptr_pop_clk_l_shift2;
	wire	[MAX_PTR_WIDTH-1:0] push_ptr_pop_clk_r_shift1;
	wire	[MAX_PTR_WIDTH-1:0] push_ptr_pop_clk_r_shift2;

	wire	[MAX_PTR_WIDTH-1:0] push_diff;
	wire	[MAX_PTR_WIDTH-1:0] push_diff_plus_1;
	wire	[MAX_PTR_WIDTH-1:0] pop_diff;
		
	wire	match_room4all;		
	wire	match_room4eight;	
	
	wire	match_one_left;			
	wire	match_one2eight_left;
	
	integer	depth_sel_push;
	integer depth_sel_pop;

  initial
  begin
    depth1_reg = DEPTH1;
    depth2_reg = DEPTH2;
    depth3_reg = DEPTH3;
  end
	
	initial
	begin
		flush_pop_clk_tf			<= 1'b0;
		push2pop_ack1					<= 1'b0;
		push2pop_ack2					<= 1'b0;
		pop_local_flush_mask	<= 1'b0;
		flush_push2pop_clk1		<= 1'b0;
		push_flush_tf_pop_clk	<= 1'b0;
		flush_push_clk_tf			<= 1'b0;
		pop2push_ack1					<= 1'b0;
		pop2push_ack2					<= 1'b0;
		push_local_flush_mask	<= 1'b0;
		flush_pop2push_clk1		<= 1'b0;
		pop_flush_tf_push_clk	<= 1'b0;
		push_ptr_push_clk			<= 0;
		pop_ptr_push_clk			<= 0;
		pop_ptr_async					<= 0;
		fifo_full_flag_f			<= 0;
		pop_ptr_pop_clk				<= 0;
		push_ptr_pop_clk			<= 0;
		push_ptr_async				<= 0;
		fifo_empty_flag_f			<= 1;
		Fifo_Full_Usr					<= 4'b0001;
		Fifo_Empty_Usr				<= 4'b0000;
	end

	assign	Fifo_Full		= fifo_full_flag_f;
	assign	Fifo_Empty	= fifo_empty_flag_f;

	assign	Write_Addr	= push_ptr_push_clk[MAX_PTR_WIDTH-2:0];
	assign	Read_Addr		= next_pop_ptr_pop_clk[MAX_PTR_WIDTH-2:0];

	assign	push_ptr_push_clk_plus1			= push_ptr_push_clk + 1;
	assign	next_push_ptr_push_clk			= ( Fifo_Push ) ? push_ptr_push_clk_plus1 : push_ptr_push_clk;
	assign	next_push_ptr_push_clk_mask	= { ( push_ptr_push_clk_mask & next_push_ptr_push_clk[MAX_PTR_WIDTH-1:MAX_PTR_WIDTH-2] ), next_push_ptr_push_clk[MAX_PTR_WIDTH-3:0] };	

	assign	pop_ptr_pop_clk_plus1				= pop_ptr_pop_clk + 1;
	assign	next_pop_ptr_pop_clk				= ( Fifo_Pop ) ? pop_ptr_pop_clk_plus1 : pop_ptr_pop_clk;
	assign	next_pop_ptr_pop_clk_mask		= { ( pop_ptr_pop_clk_mask & next_pop_ptr_pop_clk[MAX_PTR_WIDTH-1:MAX_PTR_WIDTH-2] ), next_pop_ptr_pop_clk[MAX_PTR_WIDTH-3:0] };

	assign	pop_ptr_push_clk_l_shift1	= { pop_ptr_push_clk[MAX_PTR_WIDTH-2:0], 1'b0 };
	assign	pop_ptr_push_clk_l_shift2	= { pop_ptr_push_clk[MAX_PTR_WIDTH-3:0], 2'b0 };
	assign	pop_ptr_push_clk_r_shift1	= { 1'b0, pop_ptr_push_clk[MAX_PTR_WIDTH-1:1] };
	assign	pop_ptr_push_clk_r_shift2	= { 2'b0, pop_ptr_push_clk[MAX_PTR_WIDTH-1:2] };

	assign	push_ptr_pop_clk_l_shift1	= { push_ptr_pop_clk[MAX_PTR_WIDTH-2:0], 1'b0 };
	assign	push_ptr_pop_clk_l_shift2	= { push_ptr_pop_clk[MAX_PTR_WIDTH-3:0], 2'b0 };
	assign	push_ptr_pop_clk_r_shift1	= { 1'b0, push_ptr_pop_clk[MAX_PTR_WIDTH-1:1] };
	assign	push_ptr_pop_clk_r_shift2	= { 2'b0, push_ptr_pop_clk[MAX_PTR_WIDTH-1:2] };

	assign	push_diff					= next_push_ptr_push_clk_mask - pop_ptr_push_clk_mux;
	assign	push_diff_plus_1	= push_diff + 1;
	assign	pop_diff					= push_ptr_pop_clk_mux - next_pop_ptr_pop_clk_mask;

	assign	match_room4all		= ~|push_diff;
	assign	match_room4eight	= ( depth_sel_push == 3 ) ? ( push_diff >= DEPTH3-8 ) : ( depth_sel_push == 2 ) ? ( push_diff >= DEPTH2-8 ) : ( push_diff >= DEPTH1-8 );
	
	assign	match_one_left				= ( pop_diff == 1 );
	assign	match_one2eight_left	= ( pop_diff < 8 );

	assign	push_flush_gated	= Fifo_Push_Flush & ~push_local_flush_mask;
	assign	pop_flush_gated		= Fifo_Pop_Flush & ~pop_local_flush_mask;
	
	assign	push_clk_rst	= flush_pop2push_clk1 ^ pop_flush_tf_push_clk;
	assign	pop_clk_rst		= flush_push2pop_clk1 ^ push_flush_tf_pop_clk;
	
	assign	pop_flush_done	= push2pop_ack1 ^ push2pop_ack2;
	assign	push_flush_done	= pop2push_ack1 ^ pop2push_ack2;
	
	assign	push_clk_rst_mux	= ( Fifo_Sync_Mode ) ? ( Fifo_Push_Flush | Fifo_Pop_Flush ) : ( push_flush_gated | push_clk_rst );
	assign	pop_clk_rst_mux		= ( Fifo_Sync_Mode ) ? ( Fifo_Push_Flush | Fifo_Pop_Flush ) : ( pop_flush_gated | ( pop_local_flush_mask & ~pop_flush_done ) | pop_clk_rst );
	
	//PPII
	reg match_room_at_most63, match_at_most63_left;
	
	always@( push_diff or push_diff_plus_1 or depth_sel_push or match_room4none or match_room4one )
	begin
		if( depth_sel_push == 1 ) // BR & CR: 256, DR : 512
		begin
			match_room4none		<= ( push_diff[D1_QTR_A+2:0] == depth1_reg[D1_QTR_A+2:0] );
// syao 2/12/2013
			match_room4one		<= ( push_diff_plus_1[D1_QTR_A+2:0] == depth1_reg ) | match_room4none;

			match_room4half		<= ( push_diff[D1_QTR_A+1] == 1'b1 );
			match_room4quart	<= ( push_diff[D1_QTR_A] == 1'b1 );
			//PPII
			match_room_at_most63    <=  push_diff[6];
		end
		else if( depth_sel_push == 2 ) // BR & CR : 512, DR : 1K
		begin
			match_room4none		<= ( push_diff[D2_QTR_A+2:0] == depth2_reg[D2_QTR_A+2:0] );
// syao 2/12/2013
			match_room4one		<= ( push_diff_plus_1[D2_QTR_A+2:0] == depth2_reg ) | match_room4none;

			match_room4half		<= ( push_diff[D2_QTR_A+1] == 1'b1 );
			match_room4quart	<= ( push_diff[D2_QTR_A] == 1'b1 );
			//PPII
// syao 2/12/2013
//			match_room_at_most63    <=  push_diff[6];
			match_room_at_most63    <=  &push_diff[7:6];
		end
		else  // BR & CR : 1K, DR : 2K
		begin
			match_room4none		<= ( push_diff == depth3_reg );
			match_room4one		<= ( push_diff_plus_1 == depth3_reg ) | match_room4none;

			match_room4half		<= ( push_diff[D3_QTR_A+1] == 1'b1 );
			match_room4quart	<= ( push_diff[D3_QTR_A] == 1'b1 );
			//PPII
// syao 2/12/2013
//			match_room_at_most63	<= &push_diff[7:6];
			match_room_at_most63	<= &push_diff[8:6];
		end
	end
	
	//PPII
	
	assign room4_32s = ~push_diff[5];
	assign room4_16s = ~push_diff[4];
	assign room4_8s  = ~push_diff[3];
	assign room4_4s  = ~push_diff[2];
	assign room4_2s  = ~push_diff[1];
	assign room4_1s  = &push_diff[1:0];				
	
	always@( depth_sel_pop or pop_diff )
	begin
		if( depth_sel_pop == 1 ) // BR & CR: 256, DR : 512
		begin
			match_all_left		<= ( pop_diff[D1_QTR_A+2:0] == depth1_reg[D1_QTR_A+2:0] );

			match_half_left		<= ( pop_diff[D1_QTR_A+1] == 1'b1 );
			match_quart_left	<= ( pop_diff[D1_QTR_A] == 1'b1 );
			//PPII
			match_at_most63_left	<= ~pop_diff[6];
		end
		else if( depth_sel_pop == 2 ) // BR & CR : 512, DR : 1K
		begin
			match_all_left		<= ( pop_diff[D2_QTR_A+2:0] == depth2_reg[D2_QTR_A+2:0] );

			match_half_left		<= ( pop_diff[D2_QTR_A+1] == 1'b1 );
			match_quart_left	<= ( pop_diff[D2_QTR_A] == 1'b1 );
			//PPII
// syao 2/12/2013
//			match_at_most63_left	<= ~pop_diff[6];			
			match_at_most63_left	<= ~|pop_diff[7:6];			
		end
		else  // BR & CR : 1K, DR : 2K
		begin
			match_all_left		<= ( pop_diff == depth3_reg );

			match_half_left		<= ( pop_diff[D3_QTR_A+1] == 1'b1 );
			match_quart_left	<= ( pop_diff[D3_QTR_A] == 1'b1 );
			//PPII
// syao 2/12/2013
//			match_at_most63_left	<= ~|pop_diff[7:6];			
			match_at_most63_left	<= ~|pop_diff[8:6];			
		end
	end
	
	//PPII
	
	assign at_least_32 = pop_diff[5];
	assign at_least_16 = pop_diff[4];
	assign at_least_8 = pop_diff[3];
	assign at_least_4 = pop_diff[2];
	assign at_least_2 = pop_diff[1];
	assign one_left = pop_diff[0];
	
	
	always@( posedge Pop_Clk or negedge Rst_n )
	begin
		if( ~Rst_n )
		begin
			push2pop_ack1 <= 1'b0;
			push2pop_ack2 <= 1'b0;
			flush_pop_clk_tf <= 1'b0;
			pop_local_flush_mask <= 1'b0;
			flush_push2pop_clk1 <= 1'b0;
			push_flush_tf_pop_clk <= 1'b0;
		end
		else
		begin
			push2pop_ack1 <= pop_flush_tf_push_clk;
			push2pop_ack2 <= push2pop_ack1;
			flush_push2pop_clk1 <= flush_push_clk_tf;
			if( pop_flush_gated )
			begin
				flush_pop_clk_tf	<= ~flush_pop_clk_tf;
			end
	
			if( pop_flush_gated & ~Fifo_Sync_Mode )
			begin
				pop_local_flush_mask	<= 1'b1;
			end
			else if( pop_flush_done )
			begin
				pop_local_flush_mask	<= 1'b0;
			end
	
			if( pop_clk_rst )
			begin
				push_flush_tf_pop_clk	<= ~push_flush_tf_pop_clk;
			end
		end
	end

	always@( posedge Push_Clk or negedge Rst_n )
	begin
		if( ~Rst_n )
		begin
			pop2push_ack1 <= 1'b0;
			pop2push_ack2 <= 1'b0;
			flush_push_clk_tf <= 1'b0;
			push_local_flush_mask <= 1'b0;
			flush_pop2push_clk1 <= 1'b0;
			pop_flush_tf_push_clk <= 1'b0;
		end
		else
		begin
			pop2push_ack1				<= push_flush_tf_pop_clk;
			pop2push_ack2				<= pop2push_ack1;
			flush_pop2push_clk1	<= flush_pop_clk_tf;
			if( push_flush_gated )
			begin
				flush_push_clk_tf	<= ~flush_push_clk_tf;
			end
	
			if( push_flush_gated & ~Fifo_Sync_Mode )
			begin
				push_local_flush_mask	<= 1'b1;
			end
			else if( push_flush_done )
			begin
				push_local_flush_mask	<= 1'b0;
			end
			
			if( push_clk_rst )
			begin
				pop_flush_tf_push_clk	<= ~pop_flush_tf_push_clk;
			end
		end
	end

	always@( Fifo_Push_Width or Fifo_Pop_Width or pop_ptr_push_clk_l_shift1 or pop_ptr_push_clk_l_shift2 or pop_ptr_push_clk_r_shift1 or
						pop_ptr_push_clk_r_shift2 or push_ptr_pop_clk_l_shift1 or push_ptr_pop_clk_l_shift2 or push_ptr_pop_clk_r_shift1 or push_ptr_pop_clk_r_shift2 or
						pop_ptr_push_clk or push_ptr_pop_clk )
	begin
		case( { Fifo_Push_Width, Fifo_Pop_Width } )
			4'b0001:	//	byte push halfword pop
      begin
      	push_ptr_push_clk_mask	<= 2'b11;
				pop_ptr_pop_clk_mask		<= 2'b01;
				pop_ptr_push_clk_mux		<= pop_ptr_push_clk_l_shift1;
				push_ptr_pop_clk_mux		<= push_ptr_pop_clk_r_shift1;
			end
			4'b0010:	//	byte push word pop
      begin
      	push_ptr_push_clk_mask	<= 2'b11;
				pop_ptr_pop_clk_mask		<= 2'b00;
				pop_ptr_push_clk_mux		<= pop_ptr_push_clk_l_shift2;
				push_ptr_pop_clk_mux		<= push_ptr_pop_clk_r_shift2;
			end
			4'b0100:	//	halfword push byte pop
      begin
      	push_ptr_push_clk_mask	<= 2'b01;
				pop_ptr_pop_clk_mask		<= 2'b11;
				pop_ptr_push_clk_mux		<= pop_ptr_push_clk_r_shift1;
				push_ptr_pop_clk_mux		<= push_ptr_pop_clk_l_shift1;
			end
      4'b0110:	//	halfword push word pop
      begin
      	push_ptr_push_clk_mask	<= 2'b11;
				pop_ptr_pop_clk_mask		<= 2'b01;
				pop_ptr_push_clk_mux		<= pop_ptr_push_clk_l_shift1;
				push_ptr_pop_clk_mux		<= push_ptr_pop_clk_r_shift1;
			end
			4'b1000:	//	word push byte pop
      begin
      	push_ptr_push_clk_mask	<= 2'b00;
				pop_ptr_pop_clk_mask		<= 2'b11;
				pop_ptr_push_clk_mux		<= pop_ptr_push_clk_r_shift2;
				push_ptr_pop_clk_mux		<= push_ptr_pop_clk_l_shift2;
			end
			4'b1001:	//	word push halfword pop
      begin
      	push_ptr_push_clk_mask	<= 2'b01;
				pop_ptr_pop_clk_mask		<= 2'b11;
				pop_ptr_push_clk_mux		<= pop_ptr_push_clk_r_shift1;
				push_ptr_pop_clk_mux		<= push_ptr_pop_clk_l_shift1;
			end
      default:	//	no conversion
      begin
      	push_ptr_push_clk_mask	<= 2'b11;
				pop_ptr_pop_clk_mask		<= 2'b11;
				pop_ptr_push_clk_mux		<= pop_ptr_push_clk;
				push_ptr_pop_clk_mux		<= push_ptr_pop_clk;
			end
  	endcase
	end
	
	always@( Fifo_Ram_Mode or Fifo_Push_Width )
	begin
		if( Fifo_Ram_Mode == Fifo_Push_Width[0] )
		begin
			depth_sel_push	<= 2;	// BR & CR : 512, DR : 1K
		end
		else if( Fifo_Ram_Mode == Fifo_Push_Width[1] )
		begin
			depth_sel_push	<= 1;	// BR & CR: 256, DR : 512
		end
		else
		begin
			depth_sel_push	<= 3;	// BR & CR : 1K, DR : 2K
		end
	end

	always@( Fifo_Ram_Mode or Fifo_Pop_Width )
	begin
		if( Fifo_Ram_Mode == Fifo_Pop_Width[0] )
		begin
			depth_sel_pop	<= 2;	// BR & CR : 512, DR : 1K
		end
		else if( Fifo_Ram_Mode == Fifo_Pop_Width[1] )
		begin
			depth_sel_pop	<= 1;	// BR & CR: 256, DR : 512
		end
		else
		begin
			depth_sel_pop	<= 3;	// BR & CR : 1K, DR : 2K
		end
	end

	always@( posedge Push_Clk or negedge Rst_n )
	begin
		if( ~Rst_n )
		begin
			push_ptr_push_clk	<= 0;
			pop_ptr_push_clk	<= 0;
			pop_ptr_async			<= 0;
			fifo_full_flag_f	<= 0;
		end
		else
		begin
			if( push_clk_rst_mux )
			begin
				push_ptr_push_clk	<= 0;
				pop_ptr_push_clk	<= 0;
				pop_ptr_async			<= 0;
				fifo_full_flag_f	<= 0;
			end
			else
			begin
				push_ptr_push_clk	<= next_push_ptr_push_clk; 
				pop_ptr_push_clk	<= ( Fifo_Sync_Mode ) ? next_pop_ptr_pop_clk : pop_ptr_async;
				pop_ptr_async			<= pop_ptr_pop_clk;
				fifo_full_flag_f	<= match_room4one | match_room4none;
			end
		end
	end

	always@( posedge Pop_Clk or negedge Rst_n )
	begin
		if( ~Rst_n )
		begin
			pop_ptr_pop_clk		<= 0;
			push_ptr_pop_clk	<= 0;
			push_ptr_async		<= 0;
			fifo_empty_flag_f	<= 1;
		end
		else
		begin
			if( pop_clk_rst_mux )
			begin
				pop_ptr_pop_clk		<= 0;
				push_ptr_pop_clk	<= 0;
				push_ptr_async		<= 0;
				fifo_empty_flag_f	<= 1;
			end
			else
			begin
				pop_ptr_pop_clk		<= next_pop_ptr_pop_clk;
				push_ptr_pop_clk	<= ( Fifo_Sync_Mode ) ? next_push_ptr_push_clk : push_ptr_async;
				push_ptr_async		<= push_ptr_push_clk;
				fifo_empty_flag_f	<= ( pop_diff == 1 ) | ( pop_diff == 0 );
			end
		end
	end	


	always@( posedge Push_Clk or negedge Rst_n )
	begin
		if( ~Rst_n )
		begin

			Fifo_Full_Usr	<= 4'b0001;
		end
		else
		begin
			if( match_room4none )
			begin
				Fifo_Full_Usr	<= 4'b0000;
			end
			else if( match_room4all )
			begin
				Fifo_Full_Usr	<= 4'b0001;
			end
			else if( ~match_room4half )
			begin
				Fifo_Full_Usr	<= 4'b0010;
			end
			else if( ~match_room4quart )
			begin
				Fifo_Full_Usr	<= 4'b0011;
			end
			else 
				begin
				if (match_room_at_most63)
					begin
					if (room4_32s)
						Fifo_Full_Usr <= 4'b1010;
					else if (room4_16s)
						Fifo_Full_Usr <= 4'b1011;
					else if (room4_8s)
						Fifo_Full_Usr <= 4'b1100;
					else if (room4_4s)
						Fifo_Full_Usr <= 4'b1101;
					else if (room4_2s)
						Fifo_Full_Usr <= 4'b1110;
					else if (room4_1s)
						Fifo_Full_Usr <= 4'b1111;
					else
						Fifo_Full_Usr <= 4'b1110;
					end
				else
					Fifo_Full_Usr <= 4'b0100;
				end
		end
	end


	always@( posedge Pop_Clk or negedge Rst_n )
	begin
		if( ~Rst_n )
		begin
			Fifo_Empty_Usr	<= 4'b0000;
		end
		else
		begin
			if( Fifo_Pop_Flush | ( pop_local_flush_mask & ~pop_flush_done ) | pop_clk_rst )
			begin
				Fifo_Empty_Usr	<= 4'b0000;
			end
			else 
			if( match_all_left )
			begin
				Fifo_Empty_Usr	<= 4'b1111;
			end
			else if( match_half_left )
			begin
				Fifo_Empty_Usr	<= 4'b1110;
			end
			else if( match_quart_left )
			begin
				Fifo_Empty_Usr	<= 4'b1101;
			end
			else 
				begin
				if (match_at_most63_left)
					begin
					if (at_least_32)
						Fifo_Empty_Usr	<= 4'b0110;
					else if	(at_least_16)
						Fifo_Empty_Usr	<= 4'b0101;					
					else if	(at_least_8)
						Fifo_Empty_Usr	<= 4'b0100;					
					else if	(at_least_4)
						Fifo_Empty_Usr	<= 4'b0011;					
					else if	(at_least_2)
						Fifo_Empty_Usr	<= 4'b0010;					
					else if	(one_left)
						Fifo_Empty_Usr	<= 4'b0001;
					else Fifo_Empty_Usr	<= 4'b0000;
					end
				else
					Fifo_Empty_Usr	<= 4'b1000;
				end
		end
	end
endmodule

`timescale 10 ps /1 ps

//`define ADDRWID 8
`define DATAWID 18 
`define WEWID 2
//`define DEPTH 256

module ram(
						AA,
						AB,
						CLKA,
						CLKB,
						WENA,
						WENB,
						CENA,
						CENB,
						WENBA,
						WENBB,
						DA,
						QA,
						DB,
						QB
					);


parameter ADDRWID = 8;
parameter DEPTH = (1<<ADDRWID);

	output	[`DATAWID-1:0]	QA;
	input										CLKA;
	input										CENA;
	input										WENA;
	input		[`WEWID-1:0]		WENBA;
	input		[ADDRWID-1:0]	AA;
	input		[`DATAWID-1:0]	DA;
	output	[`DATAWID-1:0]	QB;
	
	input										CLKB;
	input										CENB;
	input										WENB;
	input		[`WEWID-1:0]		WENBB;
	input		[ADDRWID-1:0]	AB;
	input		[`DATAWID-1:0]	DB;
	
	integer	i, j, k, l, m;

	wire									CEN1;
	wire									OEN1;
	wire									WEN1;
	wire	[`WEWID-1:0]		WENB1;
	wire	[ADDRWID-1:0]	A1;
	
	reg	[ADDRWID-1:0]	AddrOut1;
	wire	[`DATAWID-1:0]	I1;
	
	wire									CEN2;
	wire									OEN2;
	wire									WEN2;
	wire	[`WEWID-1:0]		WENB2;
	wire	[ADDRWID-1:0]	A2;
	
	reg	[ADDRWID-1:0]	AddrOut2;
	wire	[`DATAWID-1:0]	I2;
	
	reg		[`DATAWID-1:0]	O1, QAreg;
	reg		[`DATAWID-1:0]	O2, QBreg;
	
	reg										WEN1_f;
	reg										WEN2_f;
	reg	[ADDRWID-1:0]	A2_f;
	reg	[ADDRWID-1:0]	A1_f;
	
	wire									CEN1_SEL;
	wire									WEN1_SEL;
	wire	[ADDRWID-1:0]	A1_SEL;
	wire	[`DATAWID-1:0]	I1_SEL;
	wire	[`WEWID-1:0]		WENB1_SEL;
	
	wire									CEN2_SEL;
	wire									WEN2_SEL;
	wire	[ADDRWID-1:0]	A2_SEL;
	wire	[`DATAWID-1:0]	I2_SEL;
	wire	[`WEWID-1:0]		WENB2_SEL;
	wire  overlap;
	
	wire CLKA_d, CLKB_d, CEN1_d, CEN2_d;
	
	assign	A1_SEL    = AA;
	assign	I1_SEL    = DA;
	assign	CEN1_SEL  = CENA;
	assign	WEN1_SEL  = WENA;
	assign	WENB1_SEL = WENBA;
	
	assign	A2_SEL    = AB;
	assign	I2_SEL    = DB;
	assign	CEN2_SEL  = CENB;
	assign	WEN2_SEL  = WENB;
	assign	WENB2_SEL = WENBB;
	
	assign	CEN1	= CEN1_SEL;
	assign	OEN1	= 1'b0;                           
	assign	WEN1	= WEN1_SEL;
	assign	WENB1	= WENB1_SEL;
	assign	A1		= A1_SEL;
	assign	I1		= I1_SEL;
	
	assign	CEN2	= CEN2_SEL;
	assign	OEN2	= 1'b0;
	assign	WEN2	= WEN2_SEL;
	assign	WENB2	= WENB2_SEL;
	assign	A2		= A2_SEL;
	assign	I2		= I2_SEL;


	reg		[`DATAWID-1:0]	ram[DEPTH-1:0];
	reg		[`DATAWID-1:0]	wrData1;
	reg		[`DATAWID-1:0]	wrData2;
	wire	[`DATAWID-1:0]	tmpData1;
	wire	[`DATAWID-1:0]	tmpData2;
	
reg CENreg1, CENreg2;

assign #1 CLKA_d = CLKA;
assign #1 CLKB_d = CLKB;
// updated by sya 20130523
assign #2 CEN1_d = CEN1;
assign #2 CEN2_d = CEN2;

//PPII
assign	QA = QAreg | O1;
assign	QB = QBreg | O2;

	assign	tmpData1	= ram[A1];
	assign	tmpData2	= ram[A2];
	
	assign	overlap	= ( A1_f == A2_f ) & WEN1_f & WEN2_f;
	
	initial
	begin
		for( i = 0; i < DEPTH; i = i+1 )
		begin
			ram[i]	= 18'bxxxxxxxxxxxxxxxxxx;
		end
	end
	
	always@( WENB1 or I1 or tmpData1 )
	begin
		for( j = 0; j < 9; j = j+1 )
		begin
			wrData1[j]	<= ( WENB1[0] ) ? tmpData1[j] : I1[j];
		end
		for( l = 9; l < 19; l = l+1 )
		begin
			wrData1[l]	<= ( WENB1[1] ) ? tmpData1[l] : I1[l];
		end
	end
	
	always@( posedge CLKA )
	begin
		//O1	<= CEN1 ? 18'bxxxxxxxxxxxxxxxxxx : ram[A1];
		if( ~WEN1 & ~CEN1 )
		begin
			ram[A1]	<= wrData1[`DATAWID-1:0];
		end
	end
	
//pre-charging to 1 every clock cycle
	always@( posedge CLKA_d)
    if(~CEN1_d)
	    begin
	      O1	= 18'h3ffff;
        #100;
		    O1	= 18'h00000;
		end
	
//PPII
	always@( posedge CLKA )
		if (~CEN1)
			begin
			AddrOut1 <= A1;
			end

	always@( posedge CLKA_d)
		if (~CEN1_d)
			begin
			QAreg <= ram[AddrOut1];
			end


	always@( posedge CLKA )
	begin
		WEN1_f	<= ~WEN1 & ~CEN1;
		A1_f<= A1;
		
	end
	
	always@( WENB2 or I2 or tmpData2 )
	begin
		for( k = 0; k < 9; k = k+1 )
		begin
			wrData2[k]	<= ( WENB2[0] ) ? tmpData2[k] : I2[k];
		end
		for( m = 9; m < 19; m = m+1 )
		begin
			wrData2[m]	<= ( WENB2[1] ) ? tmpData2[m] : I2[m];
		end
	end
	
	always@( posedge CLKB )
	begin
		
		if( ~WEN2 & ~CEN2 )
		begin
			ram[A2]	<= wrData2[`DATAWID-1:0];
		end
	end

//pre-charging to 1 every clock cycle
	always@( posedge CLKB_d )
    if(~CEN2_d)
	    begin
	      O2	= 18'h3ffff;
        #100;
		    O2	= 18'h00000;
		end


//PPII
	always@( posedge CLKB )
		if (~CEN2)
			begin
			AddrOut2 <= A2;
			end

	always@( posedge CLKB_d )
		if (~CEN2_d)
			begin
			QBreg <= ram[AddrOut2];
			end

	always@( posedge CLKB )
	begin
		WEN2_f	<= ~WEN2 & ~CEN2;
		A2_f<=A2;
		
	end

	always@( A1_f or A2_f or overlap)
	begin
		if( overlap )
		begin
			ram[A1_f]	<= 18'bxxxxxxxxxxxxxxxxxx;
		end
	end

endmodule

`timescale 1 ns /10 ps
//`define ADDRWID 10
`define DATAWID 18
`define WEWID 2

module x2_model(
									Concat_En,
									
									ram0_WIDTH_SELA,
									ram0_WIDTH_SELB,
									ram0_PLRD,
									
									ram0_CEA,
									ram0_CEB,
									ram0_I,
									ram0_O,
									ram0_AA,
									ram0_AB,
									ram0_CSBA,
									ram0_CSBB,
									ram0_WENBA,
									
									ram1_WIDTH_SELA,
									ram1_WIDTH_SELB,
									ram1_PLRD,
									
									ram1_CEA,
									ram1_CEB,
									ram1_I,
									ram1_O,
									ram1_AA,
									ram1_AB,
									ram1_CSBA,
									ram1_CSBB,
									ram1_WENBA
								);

parameter ADDRWID = 10;								

	input										Concat_En;      
	
	input		[1:0]						ram0_WIDTH_SELA;
	input		[1:0]						ram0_WIDTH_SELB;
	input										ram0_PLRD;      
	input										ram0_CEA;
	input										ram0_CEB;
	input		[`DATAWID-1:0]	ram0_I;
	output	[`DATAWID-1:0]	ram0_O;
	input		[ADDRWID-1:0]	ram0_AA;
	input		[ADDRWID-1:0]	ram0_AB;
	input										ram0_CSBA;
	input										ram0_CSBB;
	input		[`WEWID-1:0]		ram0_WENBA;
	
	input		[1:0]						ram1_WIDTH_SELA;
	input		[1:0]						ram1_WIDTH_SELB;
	input										ram1_PLRD;
	input										ram1_CEA;
	input										ram1_CEB;
	input		[`DATAWID-1:0]	ram1_I;
	output	[`DATAWID-1:0]	ram1_O;
	input		[ADDRWID-1:0]	ram1_AA;
	input		[ADDRWID-1:0]	ram1_AB;
	input										ram1_CSBA;
	input										ram1_CSBB;
	input 	[`WEWID-1:0]		ram1_WENBA;
	
	reg										ram0_PLRDA_SEL;
	reg										ram0_PLRDB_SEL;
	reg										ram1_PLRDA_SEL;
	reg										ram1_PLRDB_SEL;
	reg										ram_AA_ram_SEL; 
	reg										ram_AB_ram_SEL;

	reg		[`WEWID-1:0]		ram0_WENBA_SEL;
	reg		[`WEWID-1:0]		ram0_WENBB_SEL;
	reg		[`WEWID-1:0]		ram1_WENBA_SEL;
	reg		[`WEWID-1:0]		ram1_WENBB_SEL;
	
  reg										ram0_A_x9_SEL;
  reg										ram0_B_x9_SEL;
  reg										ram1_A_x9_SEL;
  reg										ram1_B_x9_SEL;
  
	reg		[ADDRWID-3:0]	ram0_AA_SEL;
	reg		[ADDRWID-3:0]	ram0_AB_SEL;
	reg		[ADDRWID-3:0]	ram1_AA_SEL;
	reg		[ADDRWID-3:0]	ram1_AB_SEL;

	reg										ram0_AA_byte_SEL;
	reg										ram0_AB_byte_SEL;
	reg										ram1_AA_byte_SEL;
	reg										ram1_AB_byte_SEL;
	
	reg										ram0_AA_byte_SEL_Q;
	reg										ram0_AB_byte_SEL_Q;
	reg										ram1_AA_byte_SEL_Q;
	reg										ram1_AB_byte_SEL_Q;
	reg										ram0_A_mux_ctl_Q;
	reg										ram0_B_mux_ctl_Q;
	reg										ram1_A_mux_ctl_Q;
	reg										ram1_B_mux_ctl_Q;
	
  reg										ram0_O_mux_ctrl_Q;
  reg										ram1_O_mux_ctrl_Q;
  
	reg										ram_AA_ram_SEL_Q;
	reg										ram_AB_ram_SEL_Q;

	wire	[`DATAWID-1:0]	QA_1_SEL3;
	wire	[`DATAWID-1:0]	QB_0_SEL2;
	wire	[`DATAWID-1:0]	QB_1_SEL2;
  
	reg		[`DATAWID-1:0]	QA_0_Q;
	reg		[`DATAWID-1:0]	QB_0_Q;
	reg		[`DATAWID-1:0]	QA_1_Q;
	reg		[`DATAWID-1:0]	QB_1_Q;
	
	wire	[`DATAWID-1:0]	QA_0;
	wire	[`DATAWID-1:0]	QB_0;
	wire	[`DATAWID-1:0]	QA_1;
	wire	[`DATAWID-1:0]	QB_1;

	wire									ram0_CSBA_SEL;
	wire									ram0_CSBB_SEL;
	wire									ram1_CSBA_SEL;
	wire									ram1_CSBB_SEL;
	
	wire	[`DATAWID-1:0]	ram0_I_SEL1;
	wire	[`DATAWID-1:0]	ram1_I_SEL1;
	
	wire									dual_port;
	
	wire									ram0_WEBA_SEL;
	wire									ram0_WEBB_SEL;
	wire									ram1_WEBA_SEL;
	wire									ram1_WEBB_SEL;
	
	wire	[`DATAWID-1:0]	ram1_I_SEL2;
	
	wire	[`DATAWID-1:0]	QA_1_SEL2;
	wire	[`DATAWID-1:0]	QA_0_SEL1;
	wire	[`DATAWID-1:0]	QB_0_SEL1;
	wire	[`DATAWID-1:0]	QA_1_SEL1;
	wire	[`DATAWID-1:0]	QB_1_SEL1;

	wire	[`DATAWID-1:0]	QB_0_SEL3;
	wire	[`DATAWID-1:0]	QA_0_SEL2;

	initial
	begin
		QA_0_Q							<= 0;
		QB_0_Q							<= 0;
		QA_1_Q							<= 0;
		QB_1_Q							<= 0;
		ram0_AA_byte_SEL_Q	<= 0;
		ram0_A_mux_ctl_Q		<= 0;
		ram0_AB_byte_SEL_Q	<= 0;
		ram0_B_mux_ctl_Q		<= 0;
		ram1_AA_byte_SEL_Q	<= 0;
		ram1_A_mux_ctl_Q		<= 0;
		ram1_AB_byte_SEL_Q	<= 0;
		ram1_B_mux_ctl_Q		<= 0;
		ram_AA_ram_SEL_Q		<= 0;
		ram1_O_mux_ctrl_Q		<= 0;
		ram_AB_ram_SEL_Q		<= 0;
		ram0_O_mux_ctrl_Q		<= 0;
	end

	assign dual_port	= Concat_En & ~( ram0_WIDTH_SELA[1] | ram0_WIDTH_SELB[1] );
	
	assign ram0_CSBA_SEL	= ram0_CSBA;
	assign ram0_CSBB_SEL	= ram0_CSBB;
	assign ram1_CSBA_SEL	= Concat_En ? ram0_CSBA : ram1_CSBA;
	assign ram1_CSBB_SEL	= Concat_En ? ram0_CSBB : ram1_CSBB;

	assign ram0_O = QB_0_SEL3;
	assign ram1_O = dual_port ? QA_1_SEL3 : QB_1_SEL2;
	
	assign ram0_I_SEL1[8:0]		= ram0_I[8:0];
	assign ram1_I_SEL1[8:0]		= ram1_I[8:0];
	assign ram0_I_SEL1[17:9]	= ram0_AA_byte_SEL ? ram0_I[8:0] : ram0_I[17:9];
	assign ram1_I_SEL1[17:9]	= ( ( ~Concat_En & ram1_AA_byte_SEL ) | ( dual_port & ram0_AB_byte_SEL ) ) ? ram1_I[8:0] : ram1_I[17:9];
	
	assign ram1_I_SEL2	= ( Concat_En & ~ram0_WIDTH_SELA[1] ) ? ram0_I_SEL1 : ram1_I_SEL1;
	
	assign ram0_WEBA_SEL	= &ram0_WENBA_SEL;
	assign ram0_WEBB_SEL	= &ram0_WENBB_SEL;
	assign ram1_WEBA_SEL	= &ram1_WENBA_SEL;
	assign ram1_WEBB_SEL	= &ram1_WENBB_SEL;

	assign QA_0_SEL1	= ( ram0_PLRDA_SEL ) ? QA_0_Q : QA_0 ;
	assign QB_0_SEL1	= ( ram0_PLRDB_SEL ) ? QB_0_Q : QB_0 ;
	assign QA_1_SEL1	= ( ram1_PLRDA_SEL ) ? QA_1_Q : QA_1 ;
	assign QB_1_SEL1	= ( ram1_PLRDB_SEL ) ? QB_1_Q : QB_1 ;
	
  assign QA_1_SEL3	= ram1_O_mux_ctrl_Q ? QA_1_SEL2 : QA_0_SEL2;
	
	assign QA_0_SEL2[8:0]	= ram0_A_mux_ctl_Q ? QA_0_SEL1[17:9] : QA_0_SEL1[8:0] ;
	assign QB_0_SEL2[8:0]	= ram0_B_mux_ctl_Q ? QB_0_SEL1[17:9] : QB_0_SEL1[8:0] ;
	assign QA_1_SEL2[8:0]	= ram1_A_mux_ctl_Q ? QA_1_SEL1[17:9] : QA_1_SEL1[8:0] ;
	assign QB_1_SEL2[8:0]	= ram1_B_mux_ctl_Q ? QB_1_SEL1[17:9] : QB_1_SEL1[8:0] ;
	
	assign QA_0_SEL2[17:9]	= QA_0_SEL1[17:9];
	assign QB_0_SEL2[17:9]	= QB_0_SEL1[17:9];
	assign QA_1_SEL2[17:9]	= QA_1_SEL1[17:9];
	assign QB_1_SEL2[17:9]	= QB_1_SEL1[17:9];

	assign QB_0_SEL3 = ram0_O_mux_ctrl_Q ? QB_1_SEL2 : QB_0_SEL2;
	
	always@( posedge ram0_CEA )
	begin
		QA_0_Q <= QA_0;
	end
	always@( posedge ram0_CEB )
	begin
		QB_0_Q <= QB_0;
	end
	always@( posedge ram1_CEA )
	begin
		QA_1_Q <= QA_1;
	end
	always@( posedge ram1_CEB )
	begin
		QB_1_Q <= QB_1;
	end

	always@( posedge ram0_CEA )
	begin
		if( ram0_CSBA_SEL == 0 )
			ram0_AA_byte_SEL_Q	<= ram0_AA_byte_SEL;
		if( ram0_PLRDA_SEL || ( ram0_CSBA_SEL == 0 ) )
			ram0_A_mux_ctl_Q	<= ram0_A_x9_SEL & ( ram0_PLRDA_SEL ? ram0_AA_byte_SEL_Q : ram0_AA_byte_SEL );
	end
	
	always@( posedge ram0_CEB)
	begin
		if( ram0_CSBB_SEL == 0 )
			ram0_AB_byte_SEL_Q	<= ram0_AB_byte_SEL;
		if( ram0_PLRDB_SEL || ( ram0_CSBB_SEL == 0 ) )
			ram0_B_mux_ctl_Q	<= ram0_B_x9_SEL & ( ram0_PLRDB_SEL ? ram0_AB_byte_SEL_Q : ram0_AB_byte_SEL );
	end
	
	always@( posedge ram1_CEA )
	begin
		if( ram1_CSBA_SEL == 0 )
			ram1_AA_byte_SEL_Q	<= ram1_AA_byte_SEL;
		if( ram1_PLRDA_SEL || (ram1_CSBA_SEL == 0 ) )
			ram1_A_mux_ctl_Q	<= ram1_A_x9_SEL & ( ram1_PLRDA_SEL ? ram1_AA_byte_SEL_Q : ram1_AA_byte_SEL );
	end
	
	always@( posedge ram1_CEB )
	begin
		if( ram1_CSBB_SEL == 0 )
			ram1_AB_byte_SEL_Q	<= ram1_AB_byte_SEL;
		if( ram1_PLRDB_SEL || (ram1_CSBB_SEL == 0 ) )
			ram1_B_mux_ctl_Q	<= ram1_B_x9_SEL & ( ram1_PLRDB_SEL ? ram1_AB_byte_SEL_Q : ram1_AB_byte_SEL );
	end

	always@( posedge ram0_CEA )
	begin
		ram_AA_ram_SEL_Q	<= ram_AA_ram_SEL;
		ram1_O_mux_ctrl_Q	<= ( ram0_PLRDA_SEL ? ram_AA_ram_SEL_Q : ram_AA_ram_SEL );
	end

	always@( posedge ram0_CEB )
	begin
		ram_AB_ram_SEL_Q	<= ram_AB_ram_SEL;
		ram0_O_mux_ctrl_Q	<= ( ram0_PLRDB_SEL ? ram_AB_ram_SEL_Q : ram_AB_ram_SEL );
	end

	always@( Concat_En or ram0_WIDTH_SELA or ram0_WIDTH_SELB or ram0_AA or ram0_AB or ram0_WENBA or 
	         ram1_AA or ram1_AB or ram1_WENBA or ram0_PLRD or ram1_PLRD or ram1_WIDTH_SELA or ram1_WIDTH_SELB ) 
	begin
		ram0_A_x9_SEL			<= ( ~|ram0_WIDTH_SELA );
		ram1_A_x9_SEL			<= ( ~|ram0_WIDTH_SELA );
		ram0_B_x9_SEL			<= ( ~|ram0_WIDTH_SELB );
		ram0_AA_byte_SEL	<= ram0_AA[0] & ( ~|ram0_WIDTH_SELA );
		ram0_AB_byte_SEL	<= ram0_AB[0] & ( ~|ram0_WIDTH_SELB );
		if( ~Concat_En )
		begin
			ram_AA_ram_SEL	<= 1'b0;
			ram_AB_ram_SEL	<= 1'b0;
			ram1_B_x9_SEL		<= ( ~|ram1_WIDTH_SELB );
			
			ram0_PLRDA_SEL	<= ram0_PLRD;
			ram0_PLRDB_SEL	<= ram0_PLRD;
			ram1_PLRDA_SEL	<= ram1_PLRD;
			ram1_PLRDB_SEL	<= ram1_PLRD;
			ram0_WENBB_SEL	<= {`WEWID{1'b1}};
			ram1_WENBB_SEL	<= {`WEWID{1'b1}};
			
			ram0_AA_SEL				<= ram0_AA >> ( ~|ram0_WIDTH_SELA );
			ram0_WENBA_SEL[0]	<= ( ram0_AA[0] & ( ~|ram0_WIDTH_SELA ) ) | ram0_WENBA[0];
			ram0_WENBA_SEL[1]	<= ( ~ram0_AA[0] & ( ~|ram0_WIDTH_SELA ) ) | ram0_WENBA[( |ram0_WIDTH_SELA )];
			ram0_AB_SEL				<= ram0_AB >> ( ~|ram0_WIDTH_SELB );

			ram1_AA_SEL				<= ram1_AA >> ( ~|ram1_WIDTH_SELA );
			ram1_AA_byte_SEL	<= ram1_AA[0] & ( ~|ram1_WIDTH_SELA );
			ram1_WENBA_SEL[0]	<= ( ram1_AA[0] & ( ~|ram1_WIDTH_SELA ) ) | ram1_WENBA[0];
			ram1_WENBA_SEL[1]	<= ( ~ram1_AA[0] & ( ~|ram1_WIDTH_SELA ) ) | ram1_WENBA[( |ram1_WIDTH_SELA )];
			ram1_AB_SEL				<= ram1_AB >> ( ~|ram1_WIDTH_SELB );
			ram1_AB_byte_SEL	<= ram1_AB[0] & ( ~|ram1_WIDTH_SELB );
		end
		else
		begin
			ram_AA_ram_SEL	<= ~ram0_WIDTH_SELA[1] & ram0_AA[~ram0_WIDTH_SELA[0]];
			ram_AB_ram_SEL	<= ~ram0_WIDTH_SELB[1] & ram0_AB[~ram0_WIDTH_SELB[0]];
			ram1_B_x9_SEL	<= ( ~|ram0_WIDTH_SELB );

			ram0_PLRDA_SEL	<= ram1_PLRD;
			ram1_PLRDA_SEL	<= ram1_PLRD;
			ram0_PLRDB_SEL	<= ram0_PLRD;
			ram1_PLRDB_SEL	<= ram0_PLRD;
			
			ram0_AA_SEL				<= ram0_AA >> { ~ram0_WIDTH_SELA[1] & ~( ram0_WIDTH_SELA[1] ^ ram0_WIDTH_SELA[0] ), ~ram0_WIDTH_SELA[1] & ram0_WIDTH_SELA[0] };
			ram1_AA_SEL				<= ram0_AA >> { ~ram0_WIDTH_SELA[1] & ~( ram0_WIDTH_SELA[1] ^ ram0_WIDTH_SELA[0] ), ~ram0_WIDTH_SELA[1] & ram0_WIDTH_SELA[0] };
			ram1_AA_byte_SEL	<= ram0_AA[0] & ( ~|ram0_WIDTH_SELA );
			ram0_WENBA_SEL[0]	<= ram0_WENBA[0] | ( ~ram0_WIDTH_SELA[1] & ( ram0_AA[0] | ( ~ram0_WIDTH_SELA[0] & ram0_AA[1] ) ) );
			ram0_WENBA_SEL[1]	<= ( ( ~|ram0_WIDTH_SELA & ram0_WENBA[0] ) | ( |ram0_WIDTH_SELA & ram0_WENBA[1] ) ) | ( ~ram0_WIDTH_SELA[1] & ( ( ram0_WIDTH_SELA[0] & ram0_AA[0] ) | ( ~ram0_WIDTH_SELA[0] & ~ram0_AA[0] ) | ( ~ram0_WIDTH_SELA[0] & ram0_AA[1] ) ) );

			ram1_WENBA_SEL[0]	<= ( ( ~ram0_WIDTH_SELA[1] & ram0_WENBA[0] ) | ( ram0_WIDTH_SELA[1] & ram1_WENBA[0] ) ) | ( ~ram0_WIDTH_SELA[1] & ( ( ram0_WIDTH_SELA[0] & ~ram0_AA[0] ) | ( ~ram0_WIDTH_SELA[0] & ram0_AA[0] ) | ( ~ram0_WIDTH_SELA[0] & ~ram0_AA[1] ) ) );
			ram1_WENBA_SEL[1]	<= ( ( ( ram0_WIDTH_SELA == 2'b00 ) & ram0_WENBA[0] ) | ( ( ram0_WIDTH_SELA[1] == 1'b1 ) & ram1_WENBA[1] ) | ( ( ram0_WIDTH_SELA == 2'b01 ) & ram0_WENBA[1] ) ) | ( ~ram0_WIDTH_SELA[1] & ( ~ram0_AA[0] | ( ~ram0_WIDTH_SELA[0] & ~ram0_AA[1] ) ) );

			ram0_AB_SEL				<= ram0_AB >> { ~ram0_WIDTH_SELB[1] & ~( ram0_WIDTH_SELB[1] ^ ram0_WIDTH_SELB[0] ), ~ram0_WIDTH_SELB[1] & ram0_WIDTH_SELB[0] };
			ram1_AB_SEL				<= ram0_AB >> { ~ram0_WIDTH_SELB[1] & ~( ram0_WIDTH_SELB[1] ^ ram0_WIDTH_SELB[0] ), ~ram0_WIDTH_SELB[1] & ram0_WIDTH_SELB[0] };
			ram1_AB_byte_SEL	<= ram0_AB[0] & ( ~|ram0_WIDTH_SELB );
			ram0_WENBB_SEL[0]	<= ram0_WIDTH_SELB[1] | ( ram0_WIDTH_SELA[1] | ram1_WENBA[0] | ( ram0_AB[0] | ( ~ram0_WIDTH_SELB[0] & ram0_AB[1] ) ) );
			ram0_WENBB_SEL[1]	<= ram0_WIDTH_SELB[1] | ( ram0_WIDTH_SELA[1] | ( ( ~|ram0_WIDTH_SELB & ram1_WENBA[0] ) | ( |ram0_WIDTH_SELB & ram1_WENBA[1] ) ) | ( ( ram0_WIDTH_SELB[0] & ram0_AB[0] ) | ( ~ram0_WIDTH_SELB[0] & ~ram0_AB[0] ) | ( ~ram0_WIDTH_SELB[0] & ram0_AB[1] ) ) );
			ram1_WENBB_SEL[0]	<= ram0_WIDTH_SELB[1] | ( ram0_WIDTH_SELA[1] | ram1_WENBA[0] | ( ( ram0_WIDTH_SELB[0] & ~ram0_AB[0] ) | ( ~ram0_WIDTH_SELB[0] & ram0_AB[0] ) | ( ~ram0_WIDTH_SELB[0] & ~ram0_AB[1] ) ) );
			ram1_WENBB_SEL[1]	<= ram0_WIDTH_SELB[1] | ( ram0_WIDTH_SELA[1] | ( ( ~|ram0_WIDTH_SELB & ram1_WENBA[0] ) | ( |ram0_WIDTH_SELB & ram1_WENBA[1] ) ) | ( ~ram0_AB[0] | ( ~ram0_WIDTH_SELB[0] & ~ram0_AB[1] ) ) );
		end
	end
  
	

	ram	#(.ADDRWID(ADDRWID-2)) ram0_inst(
									.AA( ram0_AA_SEL ),
									.AB( ram0_AB_SEL ),
									.CLKA( ram0_CEA ),
									.CLKB( ram0_CEB ),
									.WENA( ram0_WEBA_SEL ),
									.WENB( ram0_WEBB_SEL ),
									.CENA( ram0_CSBA_SEL ),
									.CENB( ram0_CSBB_SEL ),
									.WENBA( ram0_WENBA_SEL ),
									.WENBB( ram0_WENBB_SEL ),
									.DA( ram0_I_SEL1 ),
									.QA( QA_0 ),
									.DB( ram1_I_SEL1 ),
									.QB( QB_0 )
								);

	ram	#(.ADDRWID(ADDRWID-2)) ram1_inst(
									.AA( ram1_AA_SEL ),
									.AB( ram1_AB_SEL ),
									.CLKA( ram1_CEA ),
									.CLKB( ram1_CEB ),
									.WENA( ram1_WEBA_SEL ),
									.WENB( ram1_WEBB_SEL ),
									.CENA( ram1_CSBA_SEL ),
									.CENB( ram1_CSBB_SEL ),
									.WENBA( ram1_WENBA_SEL ),
									.WENBB( ram1_WENBB_SEL ),
									.DA( ram1_I_SEL2 ),
									.QA( QA_1 ),
									.DB( ram1_I_SEL1 ),
									.QB( QB_1 )
								);


endmodule

`timescale 1 ns /10 ps
`define ADDRWID 11
`define DATAWID 18
`define WEWID 2

module ram_block_8K (  
                                CLK1_0,
                                CLK2_0,
                                WD_0,
                                RD_0,
                                A1_0,
                                A2_0,
                                CS1_0,
                                CS2_0,
                                WEN1_0,
                                POP_0,
                                Almost_Full_0,
                                Almost_Empty_0,
                                PUSH_FLAG_0,
                                POP_FLAG_0,
                                
                                FIFO_EN_0,
                                SYNC_FIFO_0,
                                PIPELINE_RD_0,
                                WIDTH_SELECT1_0,
                                WIDTH_SELECT2_0,
                                
                                CLK1_1,
                                CLK2_1,
                                WD_1,
                                RD_1,
                                A1_1,
                                A2_1,
                                CS1_1,
                                CS2_1,
                                WEN1_1,
                                POP_1,
                                Almost_Empty_1,
                                Almost_Full_1,
                                PUSH_FLAG_1,
                                POP_FLAG_1,
                                
                                FIFO_EN_1,
                                SYNC_FIFO_1,
                                PIPELINE_RD_1,
                                WIDTH_SELECT1_1,
                                WIDTH_SELECT2_1,
                                
                                CONCAT_EN_0,
                                CONCAT_EN_1,
				//PPII additional
				PUSH_0,
				PUSH_1,
				aFlushN_0,
				aFlushN_1
				
                              );

  input                   CLK1_0;
  input                   CLK2_0;
  input   [`DATAWID-1:0]  WD_0;
  output  [`DATAWID-1:0]  RD_0;
  input   [`ADDRWID-1:0]    A1_0; //chnge
  input   [`ADDRWID-1:0]    A2_0; //chnge
  input                   CS1_0;
  input                   CS2_0;
  input   [`WEWID-1:0]    WEN1_0;
  input                   POP_0;
  output                  Almost_Full_0;
  output                  Almost_Empty_0;
  output  [3:0]           PUSH_FLAG_0;
  output  [3:0]           POP_FLAG_0;
  input                   FIFO_EN_0;
  input                   SYNC_FIFO_0;
  input                   PIPELINE_RD_0;
  input   [1:0]           WIDTH_SELECT1_0;
  input   [1:0]           WIDTH_SELECT2_0;
  
  input                   CLK1_1;
  input                   CLK2_1;
  input   [`DATAWID-1:0]  WD_1;
  output  [`DATAWID-1:0]  RD_1;
  input   [`ADDRWID-1:0]    A1_1; //chnge
  input   [`ADDRWID-1:0]    A2_1; //chnge
  input                   CS1_1;
  input                   CS2_1;
  input   [`WEWID-1:0]    WEN1_1;
  input                   POP_1;
  output                  Almost_Full_1;
  output                  Almost_Empty_1;
  output  [3:0]           PUSH_FLAG_1;
  output  [3:0]           POP_FLAG_1;
  input                   FIFO_EN_1;
  input                   SYNC_FIFO_1;
  input                   PIPELINE_RD_1;
  input   [1:0]           WIDTH_SELECT1_1;
  input   [1:0]           WIDTH_SELECT2_1;
  
  input                   CONCAT_EN_0;
  input                   CONCAT_EN_1;
 
 				//PPII additional
  input                   PUSH_0;
  input                   PUSH_1;
  input                   aFlushN_0;
  input                   aFlushN_1;
  
  reg                   rstn;
    
  wire  [`WEWID-1:0]    RAM0_WENb1_SEL;
  wire  [`WEWID-1:0]    RAM1_WENb1_SEL;
  
  wire                  RAM0_CS1_SEL;
  wire                  RAM0_CS2_SEL;
  wire                  RAM1_CS1_SEL;
  wire                  RAM1_CS2_SEL;

  wire  [`ADDRWID-1:0]  Fifo0_Write_Addr;
  wire  [`ADDRWID-1:0]  Fifo0_Read_Addr;
                        
  wire  [`ADDRWID-1:0]  Fifo1_Write_Addr;
  wire  [`ADDRWID-1:0]  Fifo1_Read_Addr;

  wire  [`ADDRWID-1:0]  RAM0_AA_SEL;
  wire  [`ADDRWID-1:0]  RAM0_AB_SEL;
  wire  [`ADDRWID-1:0]  RAM1_AA_SEL;
  wire  [`ADDRWID-1:0]  RAM1_AB_SEL;
  
  wire                  Concat_En_SEL;
  
  //  To simulate POR
  initial
  begin
    rstn  = 1'b0;
    #30  rstn  = 1'b1;
  end
  
  assign fifo0_rstn = rstn & aFlushN_0;
  assign fifo1_rstn = rstn & aFlushN_1;

  assign Concat_En_SEL  = ( CONCAT_EN_0 | WIDTH_SELECT1_0[1] | WIDTH_SELECT2_0[1] )? 1'b1 : 1'b0;
  
  assign RAM0_AA_SEL  = FIFO_EN_0 ? Fifo0_Write_Addr : A1_0[`ADDRWID-1:0];
  assign RAM0_AB_SEL  = FIFO_EN_0 ? Fifo0_Read_Addr  : A2_0[`ADDRWID-1:0];
  assign RAM1_AA_SEL  = FIFO_EN_1 ? Fifo1_Write_Addr : A1_1[`ADDRWID-1:0];
  assign RAM1_AB_SEL  = FIFO_EN_1 ? Fifo1_Read_Addr  : A2_1[`ADDRWID-1:0];
  
  assign RAM0_WENb1_SEL = FIFO_EN_0 ? { `WEWID{ ~PUSH_0 } } : ~WEN1_0;
  assign RAM1_WENb1_SEL = ( FIFO_EN_1 & ~Concat_En_SEL ) ? { `WEWID{ ~PUSH_1 } } :
                          ( ( FIFO_EN_0 &  Concat_En_SEL ) ? ( WIDTH_SELECT1_0[1] ? { `WEWID{ ~PUSH_0 } } : { `WEWID{ 1'b1 } } ) : ~WEN1_1 );

  assign RAM0_CS1_SEL = ( FIFO_EN_0 ? CS1_0 : ~CS1_0 );
  assign RAM0_CS2_SEL = ( FIFO_EN_0 ? CS2_0 : ~CS2_0 );
  assign RAM1_CS1_SEL = ( FIFO_EN_1 ? CS1_1 : ~CS1_1 );
  assign RAM1_CS2_SEL = ( FIFO_EN_1 ? CS2_1 : ~CS2_1 );

  x2_model #(.ADDRWID(`ADDRWID)) x2_8K_model_inst(
                            .Concat_En( Concat_En_SEL ),
                            
                            .ram0_WIDTH_SELA( WIDTH_SELECT1_0 ),
                            .ram0_WIDTH_SELB( WIDTH_SELECT2_0 ),
                            .ram0_PLRD( PIPELINE_RD_0 ),
                            
                            .ram0_CEA( CLK1_0 ),
                            .ram0_CEB( CLK2_0 ),
                            .ram0_I( WD_0 ),
                            .ram0_O( RD_0 ),
                            .ram0_AA( RAM0_AA_SEL ),
                            .ram0_AB( RAM0_AB_SEL ),
                            .ram0_CSBA( RAM0_CS1_SEL ),
                            .ram0_CSBB( RAM0_CS2_SEL ),
                            .ram0_WENBA( RAM0_WENb1_SEL ),
                            
                            .ram1_WIDTH_SELA( WIDTH_SELECT1_1 ),
                            .ram1_WIDTH_SELB( WIDTH_SELECT2_1 ),
                            .ram1_PLRD( PIPELINE_RD_1 ),
                            
                            .ram1_CEA( CLK1_1 ),
                            .ram1_CEB( CLK2_1 ),
                            .ram1_I( WD_1 ),
                            .ram1_O( RD_1 ),
                            .ram1_AA( RAM1_AA_SEL ),
                            .ram1_AB( RAM1_AB_SEL ),
                            .ram1_CSBA( RAM1_CS1_SEL ),
                            .ram1_CSBB( RAM1_CS2_SEL ),
                            .ram1_WENBA( RAM1_WENb1_SEL )
                          );

  fifo_controller_model #(.MAX_PTR_WIDTH(`ADDRWID+1)) fifo_controller0_inst(
                                                .Push_Clk( CLK1_0 ),
                                                .Pop_Clk( CLK2_0 ),
                                                
                                                .Fifo_Push( PUSH_0 ),
                                                .Fifo_Push_Flush( CS1_0 ),
                                                .Fifo_Full( Almost_Full_0 ),
                                                .Fifo_Full_Usr( PUSH_FLAG_0 ),
                                                
                                                .Fifo_Pop( POP_0 ),
                                                .Fifo_Pop_Flush( CS2_0 ),
                                                .Fifo_Empty( Almost_Empty_0 ),
                                                .Fifo_Empty_Usr( POP_FLAG_0 ),
                                                
                                                .Write_Addr( Fifo0_Write_Addr ),
                                                
                                                .Read_Addr( Fifo0_Read_Addr ),
                                                                        
                                                .Fifo_Ram_Mode( Concat_En_SEL ),
                                                .Fifo_Sync_Mode( SYNC_FIFO_0 ),
                                                .Fifo_Push_Width( WIDTH_SELECT1_0 ),
                                                .Fifo_Pop_Width( WIDTH_SELECT2_0 ),
                                                .Rst_n( fifo0_rstn )
                                              );

  fifo_controller_model #(.MAX_PTR_WIDTH(`ADDRWID+1)) fifo_controller1_inst(
                                                .Push_Clk( CLK1_1 ),
                                                .Pop_Clk( CLK2_1 ),
                                                
                                                .Fifo_Push( PUSH_1 ),
                                                .Fifo_Push_Flush( CS1_1 ),
                                                .Fifo_Full( Almost_Full_1 ),
                                                .Fifo_Full_Usr( PUSH_FLAG_1 ),
                                                
                                                .Fifo_Pop( POP_1 ),
                                                .Fifo_Pop_Flush( CS2_1 ),
                                                .Fifo_Empty( Almost_Empty_1 ),
                                                .Fifo_Empty_Usr( POP_FLAG_1 ),
                                                
                                                .Write_Addr( Fifo1_Write_Addr ),
                                                
                                                .Read_Addr( Fifo1_Read_Addr ),
                                                                        
                                                .Fifo_Ram_Mode( 1'b0 ),
                                                .Fifo_Sync_Mode( SYNC_FIFO_1 ),
                                                .Fifo_Push_Width( { 1'b0, WIDTH_SELECT1_1[0] } ),
                                                .Fifo_Pop_Width( { 1'b0, WIDTH_SELECT2_1[0] } ),
                                                .Rst_n( fifo1_rstn )
                                              );

endmodule
//pragma synthesis_off
module sw_mux (
	port_out,
	default_port,
	alt_port,
	switch
	);
	
	output port_out;
	input default_port;
	input alt_port;
	input switch;
	
	assign port_out = switch ? alt_port : default_port;
	
endmodule
//pragma synthesis_on

`define ADDRWID_8k2 11
`define DATAWID 18
`define WEWID 2

module P_PR8K_2X1_S3B (  
        CLK1_0,
        CLK2_0,
	CLK1S_0,
        CLK2S_0,
        WD_0,
        RD_0,
        A1_0,
        A2_0,
        CS1_0,
        CS2_0,
        WEN1_0,
        CLK1EN_0,
        CLK2EN_0,
        P1_0,
        P2_0,
        Almost_Full_0,
        Almost_Empty_0,
        PUSH_FLAG_0,
        POP_FLAG_0,

        FIFO_EN_0,
        SYNC_FIFO_0,
        PIPELINE_RD_0,
        WIDTH_SELECT1_0,
        WIDTH_SELECT2_0,
        DIR_0,
        ASYNC_FLUSH_0,
	ASYNC_FLUSH_S0,

        CLK1_1,
        CLK2_1,
	CLK1S_1,
        CLK2S_1,
        WD_1,
        RD_1,
        A1_1,
        A2_1,
        CS1_1,
        CS2_1,
        WEN1_1,
        CLK1EN_1,
        CLK2EN_1,
        P1_1,
        P2_1,
        Almost_Empty_1,
        Almost_Full_1,
        PUSH_FLAG_1,
        POP_FLAG_1,

        FIFO_EN_1,
        SYNC_FIFO_1,
        PIPELINE_RD_1,
        WIDTH_SELECT1_1,
        WIDTH_SELECT2_1,
        DIR_1,
        ASYNC_FLUSH_1,
	ASYNC_FLUSH_S1,

        CONCAT_EN_0,
        CONCAT_EN_1,

		SD,
		DS,
		LS,
		SD_RB1,
		LS_RB1,
		DS_RB1,
		RMEA,
		RMEB,
		RMA,
		RMB,
		TEST1A,
		TEST1B,
		RMEA_1,
		RMEB_1,
		RMA_1,
		RMB_1,
		TEST1A_1,
		TEST1B_1
);



input                   CLK1_0;
  input                   CLK2_0;
    input                   CLK1S_0;
  input                   CLK2S_0;
  input   [`DATAWID-1:0]  WD_0;
  output  [`DATAWID-1:0]  RD_0;
  input   [`ADDRWID_8k2-1:0]  A1_0;
  input   [`ADDRWID_8k2-1:0]  A2_0;
  input                   CS1_0;
  input                   CS2_0;
  input   [`WEWID-1:0]    WEN1_0;
  input  		  CLK1EN_0;
  input                   CLK2EN_0;
  input                   P1_0;
  input                   P2_0;
  output                  Almost_Full_0;
  output                  Almost_Empty_0;
  output  [3:0]           PUSH_FLAG_0;
  output  [3:0]           POP_FLAG_0;
  input                   FIFO_EN_0;
  input                   SYNC_FIFO_0;
  input                   DIR_0;
  input                   ASYNC_FLUSH_0;
  input                   ASYNC_FLUSH_S0;
  input                   PIPELINE_RD_0;
  input   [1:0]           WIDTH_SELECT1_0;
  input   [1:0]           WIDTH_SELECT2_0;
  
  input                   CLK1_1;
  input                   CLK2_1;
  input                   CLK1S_1;
  input                   CLK2S_1;
  input   [`DATAWID-1:0]  WD_1;
  output  [`DATAWID-1:0]  RD_1;
  input   [`ADDRWID_8k2-1:0]  A1_1;
  input   [`ADDRWID_8k2-1:0]  A2_1;
  input                   CS1_1;
  input                   CS2_1;
  input   [`WEWID-1:0]    WEN1_1;
  input  		  CLK1EN_1;
  input  		  CLK2EN_1;
  input  		  P1_1;
  input  		  P2_1;
  output                  Almost_Full_1;
  output                  Almost_Empty_1;
  output  [3:0]           PUSH_FLAG_1;
  output  [3:0]           POP_FLAG_1;
  input                   FIFO_EN_1;
  input                   SYNC_FIFO_1;
  input  		  DIR_1;
  input  		  ASYNC_FLUSH_1;
  input  		  ASYNC_FLUSH_S1;
  input                   PIPELINE_RD_1;
  input   [1:0]           WIDTH_SELECT1_1;
  input   [1:0]           WIDTH_SELECT2_1;
  
  input                   CONCAT_EN_0;
  input                   CONCAT_EN_1;
  
  // New Tamar RAM Ports -- Update this once the TAMAR RAM Simulation Model is ready
  input SD,DS,LS,SD_RB1,LS_RB1,DS_RB1,RMEA,RMEB,TEST1A,TEST1B,RMEA_1,RMEB_1,TEST1A_1,TEST1B_1;
  input [3:0] RMA;
  input [3:0] RMB;
  input [3:0] RMA_1;
  input [3:0] RMB_1;
    
//pragma synthesis_off
//CODE here
reg	RAM0_domain_sw;
reg	RAM1_domain_sw;

wire CLK1P_0, CLK1P_1, CLK2P_0, CLK2P_1, ASYNC_FLUSHP_1, ASYNC_FLUSHP_0;

//**Specify block information

wire	CLK1_0_int;
wire	CLK2_0_int;
wire	CLK1S_0_int;
wire	CLK2S_0_int;
wire	CS1_0_int;
wire	CS2_0_int;
wire	CLK1EN_0_int;
wire	CLK2EN_0_int;
wire	P1_0_int;
wire	P2_0_int;
wire	FIFO_EN_0_int;
wire	SYNC_FIFO_0_int;
wire	PIPELINE_RD_0_int;
wire	WIDTH_SELECT1_0_int;
wire	WIDTH_SELECT2_0_int;
wire	DIR_0_int;
wire	ASYNC_FLUSH_0_int;
wire	ASYNC_FLUSH_S0_int;
wire	CONCAT_EN_0_int;
	
wire	CLK1_1_int;
wire	CLK2_1_int;
wire	CLK1S_1_int;
wire	CLK2S_1_int;
wire	CS1_1_int;
wire	CS2_1_int;
wire	CLK1EN_1_int;
wire	CLK2EN_1_int;
wire	P1_1_int;
wire	P2_1_int;
wire	FIFO_EN_1_int;
wire	SYNC_FIFO_1_int;
wire	PIPELINE_RD_1_int;
wire	WIDTH_SELECT1_1_int;
wire	WIDTH_SELECT2_1_int;
wire	DIR_1_int;
wire	ASYNC_FLUSH_1_int;
wire	ASYNC_FLUSH_S1_int;
wire	CONCAT_EN_1_int;

wire [17:0] WD_0_int;
wire [17:0] WD_1_int;
wire [10:0] A1_0_int;
wire [10:0] A2_0_int;
wire [10:0] A1_1_int;
wire [10:0] A2_1_int;
wire [1:0] WEN1_0_int;
wire [1:0] WEN1_1_int;


buf CLK1_0_buf( CLK1_0_int, CLK1_0);
buf CLK2_0_buf(CLK2_0_int, CLK2_0);
buf CLK1S_0_buf(CLK1S_0_int, CLK1S_0);
buf CLK2S_0_buf(CLK2S_0_int, CLK2S_0);
buf CS1_0_buf( CS1_0_int, CS1_0);
buf CS2_0_buf( CS2_0_int, CS2_0);
buf CLK1EN_0_buf(CLK1EN_0_int,CLK1EN_0);
buf CLK2EN_0_buf(CLK2EN_0_int, CLK2EN_0);
buf P1_0_buf(P1_0_int, P1_0);
buf P2_0_buf(P2_0_int, P2_0);
buf FIFO_EN_0_buf(FIFO_EN_0_int,FIFO_EN_0);
buf SYNC_FIFO_0_buf(SYNC_FIFO_0_int,SYNC_FIFO_0);
buf PIPELINE_RD_0_buf(PIPELINE_RD_0_int,PIPELINE_RD_0);
buf WIDTH_SELECT1_0_buf(WIDTH_SELECT1_0_int,WIDTH_SELECT1_0);
buf WIDTH_SELECT2_0_buf(WIDTH_SELECT2_0_int,WIDTH_SELECT2_0);
buf DIR_0_buf(DIR_0_int,DIR_0);
buf ASYNC_FLUSH_0_buf(ASYNC_FLUSH_0_int, ASYNC_FLUSH_0);
buf ASYNC_FLUSH_S0_buf(ASYNC_FLUSH_S0_int, ASYNC_FLUSH_S0);
buf CONCAT_EN_0_buf(CONCAT_EN_0_int,CONCAT_EN_0);
buf CLK1_1_buf(CLK1_1_int, CLK1_1);
buf CLK2_1_buf(CLK2_1_int,CLK2_1);
buf CLK1S_1_buf(CLK1S_1_int,CLK1S_1);
buf CLK2S_1_buf(CLK2S_1_int,CLK2S_1);
buf CS1_1_buf(CS1_1_int, CS1_1);
buf CS2_1_buf(CS2_1_int,CS2_1);
buf CLK1EN_1_buf( CLK1EN_1_int, CLK1EN_1);
buf CLK2EN_1_buf( CLK2EN_1_int,CLK2EN_1);
buf P1_1_buf(P1_1_int, P1_1);
buf P2_1_buf(P2_1_int, P2_1);
buf FIFO_EN_1_buf(FIFO_EN_1_int,FIFO_EN_1);
buf SYNC_FIFO_1_buf(SYNC_FIFO_1_int,SYNC_FIFO_1);
buf PIPELINE_RD_1_buf( PIPELINE_RD_1_int,        PIPELINE_RD_1);
buf WIDTH_SELECT1_1_buf(WIDTH_SELECT1_1_int,WIDTH_SELECT1_1);
buf WIDTH_SELECT2_1_buf(WIDTH_SELECT2_1_int,WIDTH_SELECT2_1);
buf DIR_1_buf(DIR_1_int,DIR_1);
buf ASYNC_FLUSH_1_buf(ASYNC_FLUSH_1_int,ASYNC_FLUSH_1);
buf ASYNC_FLUSH_S1_buf(ASYNC_FLUSH_S1_int,ASYNC_FLUSH_S1);
buf CONCAT_EN_1_buf(CONCAT_EN_1_int,CONCAT_EN_1);

buf WD00_buf (WD_0_int[0],WD_0[0]);
buf WD01_buf (WD_0_int[1],WD_0[1]);
buf WD02_buf (WD_0_int[2],WD_0[2]);
buf WD03_buf (WD_0_int[3],WD_0[3]);
buf WD04_buf (WD_0_int[4],WD_0[4]);
buf WD05_buf (WD_0_int[5],WD_0[5]);
buf WD06_buf (WD_0_int[6],WD_0[6]);
buf WD07_buf (WD_0_int[7],WD_0[7]);
buf WD08_buf (WD_0_int[8],WD_0[8]);
buf WD09_buf (WD_0_int[9],WD_0[9]);
buf WD011_buf (WD_0_int[11],WD_0[11]);
buf WD010_buf (WD_0_int[10],WD_0[10]);
buf WD012_buf (WD_0_int[12],WD_0[12]);
buf WD013_buf (WD_0_int[13],WD_0[13]);
buf WD014_buf (WD_0_int[14],WD_0[14]);
buf WD015_buf (WD_0_int[15],WD_0[15]);
buf WD016_buf (WD_0_int[16],WD_0[16]);
buf WD017_buf (WD_0_int[17],WD_0[17]);

buf WD10_buf (WD_1_int[0],WD_1[0]);
buf WD11_buf (WD_1_int[1],WD_1[1]);
buf WD12_buf (WD_1_int[2],WD_1[2]);
buf WD13_buf (WD_1_int[3],WD_1[3]);
buf WD14_buf (WD_1_int[4],WD_1[4]);
buf WD15_buf (WD_1_int[5],WD_1[5]);
buf WD16_buf (WD_1_int[6],WD_1[6]);
buf WD17_buf (WD_1_int[7],WD_1[7]);
buf WD18_buf (WD_1_int[8],WD_1[8]);
buf WD19_buf (WD_1_int[9],WD_1[9]);
buf WD111_buf (WD_1_int[11],WD_1[11]);
buf WD110_buf (WD_1_int[10],WD_1[10]);
buf WD112_buf (WD_1_int[12],WD_1[12]);
buf WD113_buf (WD_1_int[13],WD_1[13]);
buf WD114_buf (WD_1_int[14],WD_1[14]);
buf WD115_buf (WD_1_int[15],WD_1[15]);
buf WD116_buf (WD_1_int[16],WD_1[16]);
buf WD117_buf (WD_1_int[17],WD_1[17]);

buf A100_buf (A1_0_int[0],A1_0[0]);
buf A101_buf (A1_0_int[1],A1_0[1]);
buf A102_buf (A1_0_int[2],A1_0[2]);
buf A103_buf (A1_0_int[3],A1_0[3]);
buf A104_buf (A1_0_int[4],A1_0[4]);
buf A105_buf (A1_0_int[5],A1_0[5]);
buf A106_buf (A1_0_int[6],A1_0[6]);
buf A107_buf (A1_0_int[7],A1_0[7]);
buf A108_buf (A1_0_int[8],A1_0[8]);
buf A109_buf (A1_0_int[9],A1_0[9]);
buf A1010_buf (A1_0_int[10],A1_0[10]);

buf A110_buf (A1_1_int[0],A1_1[0]);
buf A111_buf (A1_1_int[1],A1_1[1]);
buf A112_buf (A1_1_int[2],A1_1[2]);
buf A113_buf (A1_1_int[3],A1_1[3]);
buf A114_buf (A1_1_int[4],A1_1[4]);
buf A115_buf (A1_1_int[5],A1_1[5]);
buf A116_buf (A1_1_int[6],A1_1[6]);
buf A117_buf (A1_1_int[7],A1_1[7]);
buf A118_buf (A1_1_int[8],A1_1[8]);
buf A119_buf (A1_1_int[9],A1_1[9]);
buf A1110_buf (A1_1_int[10],A1_1[10]);

buf A200_buf (A2_0_int[0],A2_0[0]);
buf A201_buf (A2_0_int[1],A2_0[1]);
buf A202_buf (A2_0_int[2],A2_0[2]);
buf A203_buf (A2_0_int[3],A2_0[3]);
buf A204_buf (A2_0_int[4],A2_0[4]);
buf A205_buf (A2_0_int[5],A2_0[5]);
buf A206_buf (A2_0_int[6],A2_0[6]);
buf A207_buf (A2_0_int[7],A2_0[7]);
buf A208_buf (A2_0_int[8],A2_0[8]);
buf A209_buf (A2_0_int[9],A2_0[9]);
buf A2010_buf (A2_0_int[10],A2_0[10]);

buf A210_buf (A2_1_int[0],A2_1[0]);
buf A211_buf (A2_1_int[1],A2_1[1]);
buf A212_buf (A2_1_int[2],A2_1[2]);
buf A213_buf (A2_1_int[3],A2_1[3]);
buf A214_buf (A2_1_int[4],A2_1[4]);
buf A215_buf (A2_1_int[5],A2_1[5]);
buf A216_buf (A2_1_int[6],A2_1[6]);
buf A217_buf (A2_1_int[7],A2_1[7]);
buf A218_buf (A2_1_int[8],A2_1[8]);
buf A219_buf (A2_1_int[9],A2_1[9]);
buf A2110_buf (A2_1_int[10],A2_1[10]);

buf WEN100_buf (WEN1_0_int[0],WEN1_0[0]);
buf WEN101_buf (WEN1_0_int[1],WEN1_0[1]);
buf WEN110_buf (WEN1_1_int[0],WEN1_1[0]);
buf WEN111_buf (WEN1_1_int[1],WEN1_1[1]);

//**************************************************************************

assign WidSel1_1 = WIDTH_SELECT1_0[1];
assign WidSel2_1 = WIDTH_SELECT2_0[1];

assign CLK1P_0 = CLK1S_0_int ? ~CLK1_0_int : CLK1_0_int;
assign CLK1P_1 = CLK1S_1_int ? ~CLK1_1_int : CLK1_1_int;
assign CLK2P_0 = CLK2S_0_int ? ~CLK2_0_int : CLK2_0_int;
assign CLK2P_1 = CLK2S_1_int ? ~CLK2_1_int : CLK2_1_int;
assign ASYNC_FLUSHP_0 = ASYNC_FLUSH_S0_int? ~ASYNC_FLUSH_0_int : ASYNC_FLUSH_0_int;
assign ASYNC_FLUSHP_1 = ASYNC_FLUSH_S1_int? ~ASYNC_FLUSH_1_int : ASYNC_FLUSH_1_int;


/* FIFO mode-only switching */
always @( CONCAT_EN_0_int or FIFO_EN_0_int or FIFO_EN_1_int or WidSel1_1 or WidSel2_1 or DIR_0_int or DIR_1_int)

begin
	if (CONCAT_EN_0_int)                                               //CONCAT enabled, only RAM0 ports are checked
		begin
		if (~FIFO_EN_0_int)                                              //RAM MODE (no switching)
			begin
			RAM0_domain_sw = 1'b0;                                           //Both Switches are on default during RAM mode
			RAM1_domain_sw = 1'b0;
			end
		else                                                               //FIFO Mode
			begin
			RAM0_domain_sw = DIR_0_int;                                       //Both Switches will get DIR_0 (primary port) during concat
			RAM1_domain_sw = DIR_0_int;
			end
		end
	else                                                                 //CONCAT disabled, RAM0 and RAM1 ports are be checked
		begin
			if (WidSel1_1 || WidSel2_1)        //AUTO-CONCAT FIFO/RAM Mode Horizontal Concatenation
				begin
				if (~FIFO_EN_0_int)                                          //RAM MODE (no switching)
					begin
					RAM0_domain_sw = 1'b0;                                       //Both Switches are on default during RAM mode
					RAM1_domain_sw = 1'b0;
					end
				else                                                           //FIFO Mode
					begin
   		 		RAM0_domain_sw = DIR_0_int;                                   //Both Switches will get DIR_0 (primary port) during concat
			  	RAM1_domain_sw = DIR_0_int;
					end
				end
			else                                                             //FIFO/RAM Individual Mode
				begin
				if (~FIFO_EN_0_int)                                          //RAM0 Mode
					RAM0_domain_sw = 1'b0;
				else                                                           //FIFO0 Mode
					RAM0_domain_sw = DIR_0_int;
				if (~FIFO_EN_1_int)                                          //RAM1 Mode
					RAM1_domain_sw = 1'b0;
				else                                                           //FIFO1 Mode
			  	RAM1_domain_sw = DIR_1_int;
				end
		end
end


assign RAM0_Clk1_gated = CLK1EN_0_int & CLK1P_0;
assign RAM0_Clk2_gated = CLK2EN_0_int & CLK2P_0;
assign RAM1_Clk1_gated = CLK1EN_1_int & CLK1P_1;
assign RAM1_Clk2_gated = CLK2EN_1_int & CLK2P_1;

//PORT1 of RAMs is designated to PUSH circuitry, while PORT2 gets POP circuitry
sw_mux RAM0_clk_sw_port1 (.port_out(RAM0_clk_port1), .default_port(RAM0_Clk1_gated), .alt_port(RAM0_Clk2_gated), .switch(RAM0_domain_sw));
sw_mux RAM0_P_sw_port1 (.port_out(RAM0_push_port1), .default_port(P1_0_int), .alt_port(P2_0_int), .switch(RAM0_domain_sw));
sw_mux RAM0_Flush_sw_port1 (.port_out(RAM0CS_Sync_Flush_port1), .default_port(CS1_0_int), .alt_port(CS2_0_int), .switch(RAM0_domain_sw));
sw_mux RAM0_WidSel0_port1 (.port_out(RAM0_Wid_Sel0_port1), .default_port(WIDTH_SELECT1_0[0]), .alt_port(WIDTH_SELECT2_0[0]), .switch(RAM0_domain_sw));
sw_mux RAM0_WidSel1_port1 (.port_out(RAM0_Wid_Sel1_port1), .default_port(WIDTH_SELECT1_0[1]), .alt_port(WIDTH_SELECT2_0[1]), .switch(RAM0_domain_sw));

sw_mux RAM0_clk_sw_port2 (.port_out(RAM0_clk_port2), .default_port(RAM0_Clk2_gated), .alt_port(RAM0_Clk1_gated), .switch(RAM0_domain_sw));
sw_mux RAM0_P_sw_port2 (.port_out(RAM0_pop_port2), .default_port(P2_0_int), .alt_port(P1_0_int), .switch(RAM0_domain_sw));
sw_mux RAM0_Flush_sw_port2 (.port_out(RAM0CS_Sync_Flush_port2), .default_port(CS2_0_int), .alt_port(CS1_0_int), .switch(RAM0_domain_sw));
sw_mux RAM0_WidSel0_port2 (.port_out(RAM0_Wid_Sel0_port2), .default_port(WIDTH_SELECT2_0[0]), .alt_port(WIDTH_SELECT1_0[0]), .switch(RAM0_domain_sw));
sw_mux RAM0_WidSel1_port2 (.port_out(RAM0_Wid_Sel1_port2), .default_port(WIDTH_SELECT2_0[1]), .alt_port(WIDTH_SELECT1_0[1]), .switch(RAM0_domain_sw));

sw_mux RAM1_clk_sw_port1 (.port_out(RAM1_clk_port1), .default_port(RAM1_Clk1_gated), .alt_port(RAM1_Clk2_gated), .switch(RAM1_domain_sw));
sw_mux RAM1_P_sw_port1 (.port_out(RAM1_push_port1), .default_port(P1_1_int), .alt_port(P2_1_int), .switch(RAM1_domain_sw));
sw_mux RAM1_Flush_sw_port1 (.port_out(RAM1CS_Sync_Flush_port1), .default_port(CS1_1_int), .alt_port(CS2_1_int), .switch(RAM1_domain_sw));
sw_mux RAM1_WidSel0_port1 (.port_out(RAM1_Wid_Sel0_port1), .default_port(WIDTH_SELECT1_1[0]), .alt_port(WIDTH_SELECT2_1[0]), .switch(RAM1_domain_sw));
sw_mux RAM1_WidSel1_port1 (.port_out(RAM1_Wid_Sel1_port1), .default_port(WIDTH_SELECT1_1[1]), .alt_port(WIDTH_SELECT2_1[1]), .switch(RAM1_domain_sw));


sw_mux RAM1_clk_sw_port2 (.port_out(RAM1_clk_port2), .default_port(RAM1_Clk2_gated), .alt_port(RAM1_Clk1_gated), .switch(RAM1_domain_sw));
sw_mux RAM1_P_sw_port2 (.port_out(RAM1_pop_port2), .default_port(P2_1_int), .alt_port(P1_1_int), .switch(RAM1_domain_sw));
sw_mux RAM1_Flush_sw_port2 (.port_out(RAM1CS_Sync_Flush_port2), .default_port(CS2_1_int), .alt_port(CS1_1_int), .switch(RAM1_domain_sw));
sw_mux RAM1_WidSel0_port2 (.port_out(RAM1_Wid_Sel0_port2), .default_port(WIDTH_SELECT2_1[0]), .alt_port(WIDTH_SELECT1_1[0]), .switch(RAM1_domain_sw));
sw_mux RAM1_WidSel1_port2 (.port_out(RAM1_Wid_Sel1_port2), .default_port(WIDTH_SELECT2_1[1]), .alt_port(WIDTH_SELECT1_1[1]), .switch(RAM1_domain_sw));



ram_block_8K ram_block_8K_inst (  
                                .CLK1_0(RAM0_clk_port1),
                                .CLK2_0(RAM0_clk_port2),
                                .WD_0(WD_0_int),
                                .RD_0(RD_0),
                                .A1_0(A1_0_int),
                                .A2_0(A2_0_int),
                                .CS1_0(RAM0CS_Sync_Flush_port1),
                                .CS2_0(RAM0CS_Sync_Flush_port2),
                                .WEN1_0(WEN1_0_int),
                                .POP_0(RAM0_pop_port2),
                                .Almost_Full_0(Almost_Full_0),
                                .Almost_Empty_0(Almost_Empty_0),
                                .PUSH_FLAG_0(PUSH_FLAG_0),
                                .POP_FLAG_0(POP_FLAG_0),
                                
                                .FIFO_EN_0(FIFO_EN_0_int),
                                .SYNC_FIFO_0(SYNC_FIFO_0_int),
                                .PIPELINE_RD_0(PIPELINE_RD_0_int),
                                .WIDTH_SELECT1_0({RAM0_Wid_Sel1_port1,RAM0_Wid_Sel0_port1}),
                                .WIDTH_SELECT2_0({RAM0_Wid_Sel1_port2,RAM0_Wid_Sel0_port2}),
                                
                                .CLK1_1(RAM1_clk_port1),
                                .CLK2_1(RAM1_clk_port2),
                                .WD_1(WD_1_int),
                                .RD_1(RD_1),
                                .A1_1(A1_1_int),
                                .A2_1(A2_1_int),
                                .CS1_1(RAM1CS_Sync_Flush_port1),
                                .CS2_1(RAM1CS_Sync_Flush_port2),
                                .WEN1_1(WEN1_1_int),
                                .POP_1(RAM1_pop_port2),
                                .Almost_Empty_1(Almost_Empty_1),
                                .Almost_Full_1(Almost_Full_1),
                                .PUSH_FLAG_1(PUSH_FLAG_1),
                                .POP_FLAG_1(POP_FLAG_1),
                                
                                .FIFO_EN_1(FIFO_EN_1_int),
                                .SYNC_FIFO_1(SYNC_FIFO_1_int),
                                .PIPELINE_RD_1(PIPELINE_RD_1_int),
                                .WIDTH_SELECT1_1({RAM1_Wid_Sel1_port1,RAM1_Wid_Sel0_port1}),
                                .WIDTH_SELECT2_1({RAM1_Wid_Sel1_port2,RAM1_Wid_Sel0_port2}),
                                
                                .CONCAT_EN_0(CONCAT_EN_0_int),
                                .CONCAT_EN_1(CONCAT_EN_1_int),
				
				//PPII additional
				.PUSH_0(RAM0_push_port1),
				.PUSH_1(RAM1_push_port1),
				.aFlushN_0(~ASYNC_FLUSHP_0),
				.aFlushN_1(~ASYNC_FLUSHP_1)
				
                              );
                              /***RAM Cell Specify Block Data***/

wire fifo0_dir1_wd_CLK2_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CLK2S_0 == 1'b1);
wire fifo0_dir1_wd_CLK2_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CLK2S_0 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b0);
wire ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b1);
wire ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b0);
wire ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b1);
wire ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b0);
wire ram01_addr1_18k_x9_vc_con_CLK1_1_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b1);
wire ram01_addr1_18k_x9_vc_con_CLK1_0_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b0);
wire ram01_addr1_18k_x9_vc_con_CLK1_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b1);
wire ram01_addr1_18k_x9_vc_con_CLK1_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b0);
wire ram01_addr1_18k_x18_vc_con_CLK1_1_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b1);
wire ram01_addr1_18k_x18_vc_con_CLK1_0_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b0);
wire ram01_addr1_18k_x18_vc_con_CLK1_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b1);
wire ram01_addr1_18k_x18_vc_con_CLK1_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b0);
wire ram0_addr1_9k_x9_no_con_CLK1_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b1);
wire ram0_addr1_9k_x9_no_con_CLK1_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b0);
wire ram01_addr1_18k_x36_hc_con_CLK1_1_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b1);
wire ram01_addr1_18k_x36_hc_con_CLK1_0_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b0);
wire ram01_addr1_18k_x36_hc_con_CLK1_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b1);
wire ram01_addr1_18k_x36_hc_con_CLK1_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_0 == 1'b0);
wire ram0_addr1_9k_x18_no_con_CLK1_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b1);
wire ram0_addr1_9k_x18_no_con_CLK1_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_0 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_0 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_0 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_0 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_0 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_0 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_0 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_0 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_0 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_0 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_0 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_0 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_1 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_1 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_0 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_0 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_0 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_0 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b0);
wire fifo0_dir0_cs_ram0_concat0_CLK2_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b1);
wire fifo0_dir0_cs_ram0_concat0_CLK2_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b0);
wire fifo0_dir0_cs_ram0_concat0_CLK1_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b1);
wire fifo0_dir0_cs_ram0_concat0_CLK1_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b0);
wire ram0_wen_CLK1_1_1 = (FIFO_EN_0 == 1'b0  && CLK1S_1 == 1'b1);
wire ram0_wen_CLK1_0_1 = (FIFO_EN_0 == 1'b0  && CLK1S_1 == 1'b0);
wire ram0_wen_CLK1_1_0 = (FIFO_EN_0 == 1'b0  && CLK1S_0 == 1'b1);
wire ram0_wen_CLK1_0_0 = (FIFO_EN_0 == 1'b0  && CLK1S_0 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_1 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_1 == 1'b0);
wire ram01_addr2_18k_x9_vc_con_CLK2_1_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b1);
wire ram01_addr2_18k_x9_vc_con_CLK2_0_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b0);
wire ram01_addr2_18k_x9_vc_con_CLK2_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b1);
wire ram01_addr2_18k_x9_vc_con_CLK2_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b0);
wire ram01_addr2_18k_x18_vc_con_CLK2_1_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b1);
wire ram01_addr2_18k_x18_vc_con_CLK2_0_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b0);
wire ram01_addr2_18k_x18_vc_con_CLK2_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b1);
wire ram01_addr2_18k_x18_vc_con_CLK2_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b0);
wire ram0_addr2_9k_x9_no_con_CLK2_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b1);
wire ram0_addr2_9k_x9_no_con_CLK2_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b0);
wire ram01_addr2_18k_x36_hc_con_CLK2_1_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b1);
wire ram01_addr2_18k_x36_hc_con_CLK2_0_1 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b0);
wire ram01_addr2_18k_x36_hc_con_CLK2_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b1);
wire ram01_addr2_18k_x36_hc_con_CLK2_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b0);
wire ram0_addr2_9k_x18_no_con_CLK2_1_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b1);
wire ram0_addr2_9k_x18_no_con_CLK2_0_0 = (FIFO_EN_0 == 1'b0  && WIDTH_SELECT2_0[1] == 1'b0 && WIDTH_SELECT2_0[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b0);
wire fifo1_dir1_wd_CLK2_1_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CLK2S_1 == 1'b1);
wire fifo1_dir1_wd_CLK2_0_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CLK2S_1 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK1S_1 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b1 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b0);
wire ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1 = (DIR_1 == 1'b0  && WIDTH_SELECT1_1[1] == 1'b0 && WIDTH_SELECT1_1[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b1);
wire ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1 = (DIR_1 == 1'b0  && WIDTH_SELECT1_1[1] == 1'b0 && WIDTH_SELECT1_1[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_1 == 1'b0);
wire ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b1);
wire ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0 = (DIR_0 == 1'b0  && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT1_0[0] == 1'b0 && CONCAT_EN_0 == 1'b1 && CLK2S_0 == 1'b0);
wire ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1 = (DIR_1 == 1'b0  && WIDTH_SELECT1_1[1] == 1'b0 && WIDTH_SELECT1_1[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b1);
wire ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1 = (DIR_1 == 1'b0  && WIDTH_SELECT1_1[1] == 1'b0 && WIDTH_SELECT1_1[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b0);
wire ram1_addr1_9k_x9_no_con_CLK1_1_1 = (FIFO_EN_1 == 1'b0  && WIDTH_SELECT1_1[1] == 1'b0 && WIDTH_SELECT1_1[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b1);
wire ram1_addr1_9k_x9_no_con_CLK1_0_1 = (FIFO_EN_1 == 1'b0  && WIDTH_SELECT1_1[1] == 1'b0 && WIDTH_SELECT1_1[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b0);
wire ram1_addr1_9k_x18_no_con_CLK1_1_1 = (FIFO_EN_1 == 1'b0  && WIDTH_SELECT1_1[1] == 1'b0 && WIDTH_SELECT1_1[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b1);
wire ram1_addr1_9k_x18_no_con_CLK1_0_1 = (FIFO_EN_1 == 1'b0  && WIDTH_SELECT1_1[1] == 1'b0 && WIDTH_SELECT1_1[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_1_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_0_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b0);
wire fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_1_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b1);
wire fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_0_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_1_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_0_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b0);
wire fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_1_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b1);
wire fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_0_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b0);
wire ram1_wen_CLK2_1_1 = (FIFO_EN_1 == 1'b0  && CLK2S_1 == 1'b1);
wire ram1_wen_CLK2_0_1 = (FIFO_EN_1 == 1'b0  && CLK2S_1 == 1'b0);
wire ram1_wen_CLK1_1_1 = (FIFO_EN_1 == 1'b0  && CLK1S_1 == 1'b1);
wire ram1_wen_CLK1_0_1 = (FIFO_EN_1 == 1'b0  && CLK1S_1 == 1'b0);
wire ram1_wen_CLK2_1_0 = (FIFO_EN_1 == 1'b0  && CLK2S_0 == 1'b1);
wire ram1_wen_CLK2_0_0 = (FIFO_EN_1 == 1'b0  && CLK2S_0 == 1'b0);
wire ram1_add2r_9k_x9_no_con_CLK2_1_1 = (FIFO_EN_1 == 1'b0  && WIDTH_SELECT2_1[1] == 1'b0 && WIDTH_SELECT2_1[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b1);
wire ram1_add2r_9k_x9_no_con_CLK2_0_1 = (FIFO_EN_1 == 1'b0  && WIDTH_SELECT2_1[1] == 1'b0 && WIDTH_SELECT2_1[0] == 1'b0 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b0);
wire ram1_addr2_9k_x18_no_con_CLK2_1_1 = (FIFO_EN_1 == 1'b0  && WIDTH_SELECT2_1[1] == 1'b0 && WIDTH_SELECT2_1[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b1);
wire ram1_addr2_9k_x18_no_con_CLK2_0_1 = (FIFO_EN_1 == 1'b0  && WIDTH_SELECT2_1[1] == 1'b0 && WIDTH_SELECT2_1[0] == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_0 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_0 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_0 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_0 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_1 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_1 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_0 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_0 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_1 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_1 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_0 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK1S_0 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat0_CLK1_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat0_CLK1_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat0_CLK1_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat0_CLK1_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_0 == 1'b0);
wire fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b1);
wire fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b0);
wire fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b1);
wire fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK1S_1 == 1'b0);
wire fifo0_dir1_p1_p2_ram1_concat0_CLK1_1_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b1);
wire fifo0_dir1_p1_p2_ram1_concat0_CLK1_0_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b0);
wire fifo0_dir0_p1_p2_ram1_concat0_CLK1_1_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b1);
wire fifo0_dir0_p1_p2_ram1_concat0_CLK1_0_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK1S_1 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_0 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_0 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_0 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_0 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_1 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_1 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_0 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_0 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_1 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_1 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_0 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && CLK2S_0 == 1'b0);
wire fifo0_dir1_p1_p2_ram0_concat0_CLK2_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b1);
wire fifo0_dir1_p1_p2_ram0_concat0_CLK2_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b0);
wire fifo0_dir0_p1_p2_ram0_concat0_CLK2_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b1);
wire fifo0_dir0_p1_p2_ram0_concat0_CLK2_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_0 == 1'b0);
wire fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_1_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b1);
wire fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_0_1 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b0);
wire fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_1_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b1);
wire fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_0_1 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[1] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b1 && CLK2S_1 == 1'b0);
wire fifo0_dir1_p1_p2_ram1_concat0_CLK2_1_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b1);
wire fifo0_dir1_p1_p2_ram1_concat0_CLK2_0_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b0);
wire fifo0_dir0_p1_p2_ram1_concat0_CLK2_1_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b1);
wire fifo0_dir0_p1_p2_ram1_concat0_CLK2_0_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && CONCAT_EN_0 == 1'b0 && CLK2S_1 == 1'b0);
wire fifo0_dir1_sync_CLK2_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && SYNC_FIFO_0 == 1'b1 && CLK2S_0 == 1'b1);
wire fifo0_dir1_sync_CLK2_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && SYNC_FIFO_0 == 1'b1 && CLK2S_0 == 1'b0);
wire fifo0_dir0_sync_CLK2_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && SYNC_FIFO_0 == 1'b1 && CLK2S_0 == 1'b1);
wire fifo0_dir0_sync_CLK2_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && SYNC_FIFO_0 == 1'b1 && CLK2S_0 == 1'b0);
wire fifo1_dir1_sync_CLK2_1_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && SYNC_FIFO_1 == 1'b1 && CLK2S_1 == 1'b1);
wire fifo1_dir1_sync_CLK2_0_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && SYNC_FIFO_1 == 1'b1 && CLK2S_1 == 1'b0);
wire fifo1_dir0_sync_CLK2_1_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && SYNC_FIFO_1 == 1'b1 && CLK2S_1 == 1'b1);
wire fifo1_dir0_sync_CLK2_0_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && SYNC_FIFO_1 == 1'b1 && CLK2S_1 == 1'b0);
wire fifo0_dir1_sync_CLK1_1_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && SYNC_FIFO_0 == 1'b1 && CLK1S_0 == 1'b1);
wire fifo0_dir1_sync_CLK1_0_0 = (DIR_0 == 1'b1  && FIFO_EN_0 == 1'b1 && SYNC_FIFO_0 == 1'b1 && CLK1S_0 == 1'b0);
wire fifo0_dir0_sync_CLK1_1_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && SYNC_FIFO_0 == 1'b1 && CLK1S_0 == 1'b1);
wire fifo0_dir0_sync_CLK1_0_0 = (DIR_0 == 1'b0  && FIFO_EN_0 == 1'b1 && SYNC_FIFO_0 == 1'b1 && CLK1S_0 == 1'b0);
wire fifo1_dir1_sync_CLK1_1_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && SYNC_FIFO_1 == 1'b1 && CLK1S_1 == 1'b1);
wire fifo1_dir1_sync_CLK1_0_1 = (DIR_1 == 1'b1  && FIFO_EN_1 == 1'b1 && SYNC_FIFO_1 == 1'b1 && CLK1S_1 == 1'b0);
wire fifo1_dir0_sync_CLK1_1_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && SYNC_FIFO_1 == 1'b1 && CLK1S_1 == 1'b1);
wire fifo1_dir0_sync_CLK1_0_1 = (DIR_1 == 1'b0  && FIFO_EN_1 == 1'b1 && SYNC_FIFO_1 == 1'b1 && CLK1S_1 == 1'b0);
specify

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[0]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[1]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[2]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[3]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[4]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[5]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[6]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[7]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[8]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[9]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[9]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[9]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[9]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[9]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[9]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[9]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[9]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[10]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[10]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[10]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[10]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[10]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[10]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[10]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[10]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[11]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[11]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[11]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[11]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[11]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[11]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[11]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[11]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[12]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[12]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[12]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[12]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[12]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[12]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[12]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[12]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[13]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[13]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[13]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[13]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[13]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[13]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[13]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[13]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[14]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[14]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[14]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[14]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[14]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[14]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[14]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[14]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[15]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[15]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[15]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[15]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[15]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[15]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[15]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[15]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[16]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[16]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[16]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[16]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[16]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[16]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[16]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[16]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[17]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[17]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[17]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[17]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[17]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => RD_1[17]) = (0,0);

if (CLK1S_0 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[17]) = (0,0);

if (CLK1S_0 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_0 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT1_0[0] == 1'b0 && WIDTH_SELECT1_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b1 && WIDTH_SELECT2_0[1] == 1'b0 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK1_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b1 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b1 && WIDTH_SELECT2_0[0] == 1'b0 && WIDTH_SELECT2_0[1] == 1'b1 && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b0  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK2S_1 == 1'b1  && CONCAT_EN_0 == 1'b0 && PIPELINE_RD_1 == 1'b0 && FIFO_EN_1 == 1'b0)
(CLK2_1 => RD_1[17]) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => Almost_Empty_1) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => Almost_Empty_1) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => Almost_Empty_1) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => Almost_Empty_1) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => POP_FLAG_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => POP_FLAG_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => POP_FLAG_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => POP_FLAG_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => POP_FLAG_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => POP_FLAG_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => POP_FLAG_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => POP_FLAG_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => POP_FLAG_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => POP_FLAG_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => POP_FLAG_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => POP_FLAG_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => POP_FLAG_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK1_1 => POP_FLAG_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => POP_FLAG_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK2_1 => POP_FLAG_1[3]) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => Almost_Full_1) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => Almost_Full_1) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => Almost_Full_1) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => Almost_Full_1) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => PUSH_FLAG_1[0]) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => PUSH_FLAG_1[0]) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => PUSH_FLAG_1[0]) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => PUSH_FLAG_1[0]) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => PUSH_FLAG_1[1]) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => PUSH_FLAG_1[1]) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => PUSH_FLAG_1[1]) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => PUSH_FLAG_1[1]) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => PUSH_FLAG_1[2]) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => PUSH_FLAG_1[2]) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => PUSH_FLAG_1[2]) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => PUSH_FLAG_1[2]) = (0,0);

if (CLK1S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => PUSH_FLAG_1[3]) = (0,0);

if (CLK1S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b0)
(CLK1_1 => PUSH_FLAG_1[3]) = (0,0);

if (CLK2S_1 == 1'b0  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => PUSH_FLAG_1[3]) = (0,0);

if (CLK2S_1 == 1'b1  && FIFO_EN_1 == 1'b1 && DIR_1 == 1'b1)
(CLK2_1 => PUSH_FLAG_1[3]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[0]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[0]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[0]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[0]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[0]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[0]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[0]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[0]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[0]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[0]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[0]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[0]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[0]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[0]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[0]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[0]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[1]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[1]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[1]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[1]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[1]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[1]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[1]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[1]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[1]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[1]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[1]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[1]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[1]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[1]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[1]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[1]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[2]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[2]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[2]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[2]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[2]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[2]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[2]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[2]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[2]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[2]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[2]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[2]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[2]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[2]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[2]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[2]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[3]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[3]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[3]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[3]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[3]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[3]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[3]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[3]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[3]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[3]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[3]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[3]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[3]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[3]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[3]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[3]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[4]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[4]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[4]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[4]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[4]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[4]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[4]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[4]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[4]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[4]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[4]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[4]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[4]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[4]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[4]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[4]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[5]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[5]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[5]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[5]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[5]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[5]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[5]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[5]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[5]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[5]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[5]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[5]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[5]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[5]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[5]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[5]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[6]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[6]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[6]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[6]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[6]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[6]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[6]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[6]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[6]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[6]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[6]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[6]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[6]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[6]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[6]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[6]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[7]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[7]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[7]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[7]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[7]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[7]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[7]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[7]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[7]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[7]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[7]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[7]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[7]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[7]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[7]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[7]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[8]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[8]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[8]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[8]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[8]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[8]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[8]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[8]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[8]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[8]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[8]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[8]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[8]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[8]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[8]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[8]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[9]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[9]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[9]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[9]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[9]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[9]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[9]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[9]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[9]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[9]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[9]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[9]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[9]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[9]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[9]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[9]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[10]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[10]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[10]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[10]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[10]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[10]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[10]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[10]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[10]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[10]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[10]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[10]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[10]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[10]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[10]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[10]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[11]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[11]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[11]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[11]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[11]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[11]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[11]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[11]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[11]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[11]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[11]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[11]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[11]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[11]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[11]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[11]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[12]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[12]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[12]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[12]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[12]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[12]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[12]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[12]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[12]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[12]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[12]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[12]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[12]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[12]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[12]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[12]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[13]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[13]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[13]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[13]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[13]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[13]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[13]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[13]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[13]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[13]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[13]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[13]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[13]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[13]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[13]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[13]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[14]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[14]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[14]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[14]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[14]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[14]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[14]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[14]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[14]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[14]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[14]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[14]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[14]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[14]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[14]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[14]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[15]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[15]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[15]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[15]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[15]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[15]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[15]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[15]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[15]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[15]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[15]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[15]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[15]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[15]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[15]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[15]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[16]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[16]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[16]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[16]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[16]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[16]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[16]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[16]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[16]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[16]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[16]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[16]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[16]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[16]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[16]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[16]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[17]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[17]) = (0,0);

if (CLK1S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[17]) = (0,0);

if (CLK1S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => RD_0[17]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[17]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[17]) = (0,0);

if (CLK1S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[17]) = (0,0);

if (CLK1S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_1 => RD_0[17]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[17]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[17]) = (0,0);

if (CLK2S_0 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[17]) = (0,0);

if (CLK2S_0 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_0 => RD_0[17]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[17]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[17]) = (0,0);

if (CLK2S_1 == 1'b0  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[17]) = (0,0);

if (CLK2S_1 == 1'b1  && PIPELINE_RD_0 == 1'b0 && DIR_0 == 1'b0)
(CLK2_1 => RD_0[17]) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => Almost_Empty_0) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => Almost_Empty_0) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => Almost_Empty_0) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => Almost_Empty_0) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => POP_FLAG_0[0]) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => POP_FLAG_0[0]) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => POP_FLAG_0[0]) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => POP_FLAG_0[0]) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => POP_FLAG_0[1]) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => POP_FLAG_0[1]) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => POP_FLAG_0[1]) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => POP_FLAG_0[1]) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => POP_FLAG_0[2]) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => POP_FLAG_0[2]) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => POP_FLAG_0[2]) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => POP_FLAG_0[2]) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => POP_FLAG_0[3]) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK1_0 => POP_FLAG_0[3]) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => POP_FLAG_0[3]) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK2_0 => POP_FLAG_0[3]) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => Almost_Full_0) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => Almost_Full_0) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => Almost_Full_0) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => Almost_Full_0) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => PUSH_FLAG_0[0]) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => PUSH_FLAG_0[0]) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => PUSH_FLAG_0[0]) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => PUSH_FLAG_0[0]) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => PUSH_FLAG_0[1]) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => PUSH_FLAG_0[1]) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => PUSH_FLAG_0[1]) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => PUSH_FLAG_0[1]) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => PUSH_FLAG_0[2]) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => PUSH_FLAG_0[2]) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => PUSH_FLAG_0[2]) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => PUSH_FLAG_0[2]) = (0,0);

if (CLK1S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => PUSH_FLAG_0[3]) = (0,0);

if (CLK1S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b0)
(CLK1_0 => PUSH_FLAG_0[3]) = (0,0);

if (CLK2S_0 == 1'b0  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => PUSH_FLAG_0[3]) = (0,0);

if (CLK2S_0 == 1'b1  && FIFO_EN_0 == 1'b1 && DIR_0 == 1'b1)
(CLK2_0 => PUSH_FLAG_0[3]) = (0,0);

$hold( negedge CLK2_0, posedge WD_0[17] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[17] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[17] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[17] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[17], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[17], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[17], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[17], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[17], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[17], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[17], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[17], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[17], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[17], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[17], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[17], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[17], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[17], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[17], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[17], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[17] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[17] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[17] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[17] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[17], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[17], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[17], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[17], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[16] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[16] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[16] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[16] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[16], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[16], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[16], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[16], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[16], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[16], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[16], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[16], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[16], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[16], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[16], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[16], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[16], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[16], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[16], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[16], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[16] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[16] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[16] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[16] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[16], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[16], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[16], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[16], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[15] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[15] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[15] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[15] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[15], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[15], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[15], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[15], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[15], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[15], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[15], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[15], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[15], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[15], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[15], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[15], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[15], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[15], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[15], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[15], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[15] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[15] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[15] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[15] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[15], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[15], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[15], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[15], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[14] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[14] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[14] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[14] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[14], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[14], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[14], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[14], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[14], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[14], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[14], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[14], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[14], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[14], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[14], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[14], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[14], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[14], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[14], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[14], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[14] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[14] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[14] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[14] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[14], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[14], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[14], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[14], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[13] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[13] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[13] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[13] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[13], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[13], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[13], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[13], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[13], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[13], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[13], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[13], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[13], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[13], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[13], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[13], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[13], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[13], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[13], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[13], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[13] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[13] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[13] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[13] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[13], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[13], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[13], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[13], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[12] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[12] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[12] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[12] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[12], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[12], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[12], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[12], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[12], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[12], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[12], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[12], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[12], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[12], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[12], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[12], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[12], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[12], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[12], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[12], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[12] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[12] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[12] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[12] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[12], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[12], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[12], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[12], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[11] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[11] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[11] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[11] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[11], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[11], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[11], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[11], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[11], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[11], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[11], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[11], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[11], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[11], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[11], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[11], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[11], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[11], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[11], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[11], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[11] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[11] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[11] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[11] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[11], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[11], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[11], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[11], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[10] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[10] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[10] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[10] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[10], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[10], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[10], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[10], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[10], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[10], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[10], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[10], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[10], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[10], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[10], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[10], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[10], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[10], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[10], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[10], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[10] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[10] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[10] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[10] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[10], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[10], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[10], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[10], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[9] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[9] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[9] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[9] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[9], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[9], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[9], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[9], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[9], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[9], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[9], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[9], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[9], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[9], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[9], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[9], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[9], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[9], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[9], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[9], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[9] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[9] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[9] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[9] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[9], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[9], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[9], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[9], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[8] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[8] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[8] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[8] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[8], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[8], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[8], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[8], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[8], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[8], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[8], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[8], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[8], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[8], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[8], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[8], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[8] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[8] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[8], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[8], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[7] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[7] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[7] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[7] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[7], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[7], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[7], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[7], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[7], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[7], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[7], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[7], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[7], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[7], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[7], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[7], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[7] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[7] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[7], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[7], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[6] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[6] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[6] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[6] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[6], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[6], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[6], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[6], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[6], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[6], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[6], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[6], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[6], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[6], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[6], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[6], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[6] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[6] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[6], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[6], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[5] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[5] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[5] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[5] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[5], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[5], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[5], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[5], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[5], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[5], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[5], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[5], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[5], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[5], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[5], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[5], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[5] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[5] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[5], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[5], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[4] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[4] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[4] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[4] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[4], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[4], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[4], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[4], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[4], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[4], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[4], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[4], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[4], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[4], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[4], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[4], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[4] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[4] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[4], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[4], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[3] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[3] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[3] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[3] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[3], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[3], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[3], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[3], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[3], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[3], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[3], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[3], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[3], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[3], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[3], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[3], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[3] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[3] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[3], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[3], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[2] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[2] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[2] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[2] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[2], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[2], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[2], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[2], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[2], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[2], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[2], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[2], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[2], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[2], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[2], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[2], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[2] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[2] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[2], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[2], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[1] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[1] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[1] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[1] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[1], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[1], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[1], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[1], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[1], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[1], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[1], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[1], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[1], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[1], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[1], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[1], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[1] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[1] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[1], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[1], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge WD_0[0] &&& fifo0_dir1_wd_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_0[0] &&& fifo0_dir1_wd_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_0[0] &&& fifo0_dir1_wd_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_0[0] &&& fifo0_dir1_wd_CLK2_0_0, 0);


$setup( posedge WD_0[0], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);
$setup( negedge WD_0[0], negedge CLK2_0 &&& fifo0_dir1_wd_CLK2_1_0, 0);


$setup( posedge WD_0[0], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);
$setup( negedge WD_0[0], posedge CLK2_0 &&& fifo0_dir1_wd_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[0], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[0], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[0], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[0], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge WD_0[0], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge WD_0[0], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge WD_0[0], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge WD_0[0], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WD_0[0] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WD_0[0] &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge WD_0[0], negedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge WD_0[0], posedge CLK1_0 &&& ram0_fifo_dir0_wd_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[10] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[10] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[10] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[10] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[10], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[10], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[10], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[10], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[10] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[10] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[10] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[10] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[10], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[10], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[10], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[10], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[9] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[9] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[9] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[9] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[9], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[9], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[9], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[9], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[9] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[9] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[9] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[9] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[9], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[9], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[9], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[9], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[9] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[9] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[9] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[9] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[9], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[9], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[9], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[9], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[9] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[9] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[9] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[9] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[9], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[9], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[9], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[9], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[9] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[9] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[9] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[9] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[9], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[9], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[9], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[9], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[8] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[8] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[8] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[8] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge A1_0[8], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge A1_0[8], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge A1_0[8], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge A1_0[8], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[8] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[8] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[8] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[8] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge A1_0[8], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge A1_0[8], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge A1_0[8], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge A1_0[8], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[8] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[8] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[8] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[8] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[8], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[8], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[8], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[8], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[8] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[8] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[8] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[8] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[8], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[8], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[8], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[8], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[8] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[8] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[8] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[8] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[8], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[8], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[8], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[8], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[8] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[8] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[8] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[8] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[8], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[8], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[8], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[8], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[8] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[8] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[8] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[8] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[8], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[8], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[8], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[8], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[8] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[8] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[8] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[8] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[8], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[8], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[8], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[8], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[7] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[7] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[7] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[7] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge A1_0[7], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge A1_0[7], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge A1_0[7], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge A1_0[7], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[7] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[7] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[7] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[7] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge A1_0[7], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge A1_0[7], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge A1_0[7], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge A1_0[7], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[7] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[7] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[7] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[7] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[7], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[7], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[7], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[7], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[7] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[7] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[7] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[7] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[7], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[7], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[7], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[7], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[7] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[7] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[7] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[7] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[7], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[7], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[7], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[7], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[7] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[7] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[7] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[7] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[7], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[7], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[7], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[7], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[7] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[7] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[7] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[7] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[7], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[7], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[7], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[7], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[7] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[7] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[7] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[7] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[7], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[7], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[7], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[7], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[6] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[6] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[6] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[6] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge A1_0[6], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge A1_0[6], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge A1_0[6], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge A1_0[6], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[6] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[6] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[6] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[6] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge A1_0[6], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge A1_0[6], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge A1_0[6], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge A1_0[6], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[6] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[6] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[6] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[6] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[6], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[6], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[6], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[6], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[6] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[6] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[6] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[6] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[6], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[6], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[6], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[6], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[6] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[6] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[6] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[6] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[6], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[6], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[6], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[6], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[6] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[6] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[6] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[6] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[6], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[6], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[6], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[6], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[6] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[6] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[6] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[6] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[6], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[6], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[6], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[6], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[6] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[6] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[6] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[6] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[6], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[6], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[6], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[6], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[5] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[5] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[5] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[5] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge A1_0[5], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge A1_0[5], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge A1_0[5], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge A1_0[5], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[5] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[5] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[5] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[5] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge A1_0[5], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge A1_0[5], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge A1_0[5], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge A1_0[5], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[5] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[5] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[5] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[5] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[5], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[5], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[5], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[5], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[5] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[5] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[5] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[5] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[5], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[5], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[5], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[5], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[5] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[5] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[5] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[5] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[5], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[5], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[5], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[5], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[5] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[5] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[5] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[5] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[5], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[5], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[5], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[5], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[5] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[5] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[5] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[5] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[5], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[5], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[5], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[5], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[5] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[5] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[5] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[5] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[5], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[5], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[5], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[5], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[4] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[4] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[4] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[4] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge A1_0[4], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge A1_0[4], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge A1_0[4], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge A1_0[4], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[4] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[4] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[4] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[4] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge A1_0[4], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge A1_0[4], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge A1_0[4], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge A1_0[4], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[4] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[4] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[4] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[4] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[4], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[4], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[4], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[4], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[4] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[4] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[4] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[4] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[4], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[4], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[4], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[4], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[4] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[4] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[4] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[4] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[4], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[4], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[4], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[4], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[4] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[4] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[4] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[4] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[4], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[4], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[4], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[4], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[4] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[4] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[4] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[4] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[4], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[4], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[4], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[4], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[4] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[4] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[4] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[4] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[4], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[4], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[4], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[4], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[3] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[3] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[3] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[3] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge A1_0[3], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge A1_0[3], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge A1_0[3], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge A1_0[3], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[3] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[3] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[3] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[3] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge A1_0[3], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge A1_0[3], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge A1_0[3], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge A1_0[3], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[3] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[3] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[3] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[3] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[3], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[3], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[3], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[3], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[3] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[3] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[3] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[3] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[3], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[3], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[3], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[3], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[3] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[3] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[3] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[3] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[3], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[3], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[3], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[3], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[3] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[3] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[3] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[3] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[3], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[3], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[3], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[3], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[3] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[3] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[3] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[3] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[3], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[3], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[3], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[3], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[3] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[3] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[3] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[3] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[3], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[3], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[3], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[3], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[2] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[2] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[2] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[2] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge A1_0[2], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge A1_0[2], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge A1_0[2], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge A1_0[2], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[2] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[2] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[2] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[2] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge A1_0[2], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge A1_0[2], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge A1_0[2], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge A1_0[2], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[2] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[2] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[2] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[2] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[2], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[2], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[2], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[2], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[2] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[2] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[2] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[2] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[2], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[2], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[2], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[2], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[2] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[2] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[2] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[2] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[2], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[2], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[2], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[2], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[2] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[2] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[2] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[2] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[2], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[2], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[2], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[2], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[2] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[2] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[2] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[2] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[2], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[2], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[2], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[2], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[2] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[2] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[2] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[2] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[2], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[2], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[2], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[2], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[1] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[1] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[1] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[1] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge A1_0[1], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge A1_0[1], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge A1_0[1], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge A1_0[1], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[1] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[1] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[1] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[1] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge A1_0[1], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge A1_0[1], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge A1_0[1], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge A1_0[1], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[1] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[1] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[1] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[1] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[1], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[1], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[1], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[1], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[1] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[1] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[1] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[1] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[1], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[1], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[1], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[1], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[1] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[1] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[1] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[1] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[1], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[1], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[1], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[1], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[1] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[1] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[1] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[1] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[1], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[1], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[1], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[1], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[1] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[1] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[1] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[1] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[1], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[1], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[1], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[1], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[1] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[1] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[1] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[1] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[1], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[1], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[1], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[1], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[0] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[0] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[0] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[0] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge A1_0[0], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge A1_0[0], negedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge A1_0[0], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge A1_0[0], posedge CLK1_1 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[0] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[0] &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[0] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[0] &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$setup( posedge A1_0[0], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);
$setup( negedge A1_0[0], negedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_1_0, 0);


$setup( posedge A1_0[0], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);
$setup( negedge A1_0[0], posedge CLK1_0 &&& ram01_addr1_18k_x36_hc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[0] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[0] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[0] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[0] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[0], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[0], negedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[0], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[0], posedge CLK1_1 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[0] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[0] &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[0] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[0] &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[0], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[0], negedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[0], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[0], posedge CLK1_0 &&& ram01_addr1_18k_x18_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge A1_0[0] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_0[0] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_0[0] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_0[0] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$setup( posedge A1_0[0], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);
$setup( negedge A1_0[0], negedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_1, 0);


$setup( posedge A1_0[0], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);
$setup( negedge A1_0[0], posedge CLK1_1 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge A1_0[0] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[0] &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[0] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[0] &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$setup( posedge A1_0[0], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);
$setup( negedge A1_0[0], negedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_1_0, 0);


$setup( posedge A1_0[0], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);
$setup( negedge A1_0[0], posedge CLK1_0 &&& ram01_addr1_18k_x9_vc_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[0] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[0] &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[0] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[0] &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[0], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[0], negedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[0], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[0], posedge CLK1_0 &&& ram0_addr1_9k_x18_no_con_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge A1_0[0] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge A1_0[0] &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge A1_0[0] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge A1_0[0] &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$setup( posedge A1_0[0], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);
$setup( negedge A1_0[0], negedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_1_0, 0);


$setup( posedge A1_0[0], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);
$setup( negedge A1_0[0], posedge CLK1_0 &&& ram0_addr1_9k_x9_no_con_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);


$setup( posedge CS1_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);
$setup( negedge CS1_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);


$setup( posedge CS1_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);
$setup( negedge CS1_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);


$setup( posedge CS1_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);
$setup( negedge CS1_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);


$setup( posedge CS1_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);
$setup( negedge CS1_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);


$hold( negedge CLK2_1, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_1, 0);


$setup( posedge CS1_0, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_1, 0);
$setup( negedge CS1_0, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_1, 0);


$setup( posedge CS1_0, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_1, 0);
$setup( negedge CS1_0, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);


$setup( posedge CS1_0, negedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);
$setup( negedge CS1_0, negedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);


$setup( posedge CS1_0, posedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);
$setup( negedge CS1_0, posedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);


$setup( posedge CS1_0, negedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);
$setup( negedge CS1_0, negedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);


$setup( posedge CS1_0, posedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);
$setup( negedge CS1_0, posedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);


$setup( posedge CS1_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);
$setup( negedge CS1_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);


$setup( posedge CS1_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);
$setup( negedge CS1_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);


$setup( posedge CS1_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);
$setup( negedge CS1_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);


$setup( posedge CS1_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);
$setup( negedge CS1_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);


$hold( negedge CLK2_1, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_1, 0);


$setup( posedge CS1_0, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_1, 0);
$setup( negedge CS1_0, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_1, 0);


$setup( posedge CS1_0, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_1, 0);
$setup( negedge CS1_0, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);


$setup( posedge CS1_0, negedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);
$setup( negedge CS1_0, negedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);


$setup( posedge CS1_0, posedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);
$setup( negedge CS1_0, posedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);


$setup( posedge CS1_0, negedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);
$setup( negedge CS1_0, negedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);


$setup( posedge CS1_0, posedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);
$setup( negedge CS1_0, posedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_0_0, 0);


$setup( posedge CS1_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_1_0, 0);
$setup( negedge CS1_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_1_0, 0);


$setup( posedge CS1_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_0_0, 0);
$setup( negedge CS1_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_0_0, 0);


$setup( posedge CS1_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_1_0, 0);
$setup( negedge CS1_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_1_0, 0);


$setup( posedge CS1_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_0_0, 0);
$setup( negedge CS1_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge CS1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_0_0, 0);


$setup( posedge CS1_0, negedge CLK2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_1_0, 0);
$setup( negedge CS1_0, negedge CLK2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_1_0, 0);


$setup( posedge CS1_0, posedge CLK2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_0_0, 0);
$setup( negedge CS1_0, posedge CLK2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_0_0, 0);


$setup( posedge CS1_0, negedge CLK1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_1_0, 0);
$setup( negedge CS1_0, negedge CLK1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_1_0, 0);


$setup( posedge CS1_0, posedge CLK1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_0_0, 0);
$setup( negedge CS1_0, posedge CLK1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WEN1_0[1] &&& ram0_wen_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WEN1_0[1] &&& ram0_wen_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WEN1_0[1] &&& ram0_wen_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WEN1_0[1] &&& ram0_wen_CLK1_0_1, 0);


$setup( posedge WEN1_0[1], negedge CLK1_1 &&& ram0_wen_CLK1_1_1, 0);
$setup( negedge WEN1_0[1], negedge CLK1_1 &&& ram0_wen_CLK1_1_1, 0);


$setup( posedge WEN1_0[1], posedge CLK1_1 &&& ram0_wen_CLK1_0_1, 0);
$setup( negedge WEN1_0[1], posedge CLK1_1 &&& ram0_wen_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WEN1_0[1] &&& ram0_wen_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WEN1_0[1] &&& ram0_wen_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WEN1_0[1] &&& ram0_wen_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WEN1_0[1] &&& ram0_wen_CLK1_0_0, 0);


$setup( posedge WEN1_0[1], negedge CLK1_0 &&& ram0_wen_CLK1_1_0, 0);
$setup( negedge WEN1_0[1], negedge CLK1_0 &&& ram0_wen_CLK1_1_0, 0);


$setup( posedge WEN1_0[1], posedge CLK1_0 &&& ram0_wen_CLK1_0_0, 0);
$setup( negedge WEN1_0[1], posedge CLK1_0 &&& ram0_wen_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge WEN1_0[0] &&& ram0_wen_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WEN1_0[0] &&& ram0_wen_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WEN1_0[0] &&& ram0_wen_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WEN1_0[0] &&& ram0_wen_CLK1_0_1, 0);


$setup( posedge WEN1_0[0], negedge CLK1_1 &&& ram0_wen_CLK1_1_1, 0);
$setup( negedge WEN1_0[0], negedge CLK1_1 &&& ram0_wen_CLK1_1_1, 0);


$setup( posedge WEN1_0[0], posedge CLK1_1 &&& ram0_wen_CLK1_0_1, 0);
$setup( negedge WEN1_0[0], posedge CLK1_1 &&& ram0_wen_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge WEN1_0[0] &&& ram0_wen_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge WEN1_0[0] &&& ram0_wen_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge WEN1_0[0] &&& ram0_wen_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge WEN1_0[0] &&& ram0_wen_CLK1_0_0, 0);


$setup( posedge WEN1_0[0], negedge CLK1_0 &&& ram0_wen_CLK1_1_0, 0);
$setup( negedge WEN1_0[0], negedge CLK1_0 &&& ram0_wen_CLK1_1_0, 0);


$setup( posedge WEN1_0[0], posedge CLK1_0 &&& ram0_wen_CLK1_0_0, 0);
$setup( negedge WEN1_0[0], posedge CLK1_0 &&& ram0_wen_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_1, 0);


$setup( posedge CS2_0, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_1, 0);
$setup( negedge CS2_0, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_1, 0);


$setup( posedge CS2_0, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_1, 0);
$setup( negedge CS2_0, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_1, 0);


$hold( negedge CLK2_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);


$setup( posedge CS2_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);
$setup( negedge CS2_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);


$setup( posedge CS2_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);
$setup( negedge CS2_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);


$setup( posedge CS2_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);
$setup( negedge CS2_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);


$setup( posedge CS2_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);
$setup( negedge CS2_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);


$setup( posedge CS2_0, negedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);
$setup( negedge CS2_0, negedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_1_0, 0);


$setup( posedge CS2_0, posedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);
$setup( negedge CS2_0, posedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);


$setup( posedge CS2_0, negedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);
$setup( negedge CS2_0, negedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_1_0, 0);


$setup( posedge CS2_0, posedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);
$setup( negedge CS2_0, posedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_hc_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_1, 0);


$setup( posedge CS2_0, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_1, 0);
$setup( negedge CS2_0, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_1, 0);


$setup( posedge CS2_0, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_1, 0);
$setup( negedge CS2_0, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_1, 0);


$hold( negedge CLK2_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);


$setup( posedge CS2_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);
$setup( negedge CS2_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);


$setup( posedge CS2_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);
$setup( negedge CS2_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);


$setup( posedge CS2_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);
$setup( negedge CS2_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);


$setup( posedge CS2_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);
$setup( negedge CS2_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);


$setup( posedge CS2_0, negedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);
$setup( negedge CS2_0, negedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_1_0, 0);


$setup( posedge CS2_0, posedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);
$setup( negedge CS2_0, posedge CLK2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS2_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);


$setup( posedge CS2_0, negedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);
$setup( negedge CS2_0, negedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_1_0, 0);


$setup( posedge CS2_0, posedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);
$setup( negedge CS2_0, posedge CLK1_0 &&& fifo0_dir0_cs1_cs2_ram0_concat1_vc_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_0_0, 0);


$setup( posedge CS2_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_1_0, 0);
$setup( negedge CS2_0, negedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_1_0, 0);


$setup( posedge CS2_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_0_0, 0);
$setup( negedge CS2_0, posedge CLK2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS2_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_0_0, 0);


$setup( posedge CS2_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_1_0, 0);
$setup( negedge CS2_0, negedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_1_0, 0);


$setup( posedge CS2_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_0_0, 0);
$setup( negedge CS2_0, posedge CLK1_0 &&& fifo0_dir1_cs1_cs2_ram0_concat0_CLK1_0_0, 0);


$hold( negedge CLK2_0, posedge CS2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge CS2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge CS2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge CS2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_0_0, 0);


$setup( posedge CS2_0, negedge CLK2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_1_0, 0);
$setup( negedge CS2_0, negedge CLK2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_1_0, 0);


$setup( posedge CS2_0, posedge CLK2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_0_0, 0);
$setup( negedge CS2_0, posedge CLK2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK2_0_0, 0);


$hold( negedge CLK1_0, posedge CS2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge CS2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge CS2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge CS2_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_0_0, 0);


$setup( posedge CS2_0, negedge CLK1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_1_0, 0);
$setup( negedge CS2_0, negedge CLK1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_1_0, 0);


$setup( posedge CS2_0, posedge CLK1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_0_0, 0);
$setup( negedge CS2_0, posedge CLK1_0 &&& fifo0_dir0_cs_ram0_concat0_CLK1_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[10] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[10] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[10] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[10] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[10], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[10], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[10], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[10], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[10] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[10] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[10] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[10] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[10], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[10], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[10], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[10], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[9] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[9] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[9] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[9] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[9], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[9], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[9], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[9], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[9] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[9] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[9] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[9] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[9], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[9], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[9], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[9], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[9] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[9] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[9] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[9] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[9], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[9], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[9], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[9], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[9] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[9] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[9] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[9] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[9], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[9], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[9], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[9], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[9] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[9] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[9] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[9] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[9], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[9], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[9], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[9], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[8] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[8] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[8] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[8] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$setup( posedge A2_0[8], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$setup( negedge A2_0[8], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$setup( posedge A2_0[8], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$setup( negedge A2_0[8], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[8] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[8] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[8] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[8] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$setup( posedge A2_0[8], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$setup( negedge A2_0[8], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$setup( posedge A2_0[8], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$setup( negedge A2_0[8], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[8] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[8] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[8] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[8] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[8], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[8], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[8], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[8], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[8] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[8] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[8] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[8] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[8], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[8], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[8], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[8], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[8] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[8] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[8] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[8] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[8], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[8], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[8], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[8], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[8] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[8] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[8] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[8] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[8], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[8], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[8], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[8], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[8] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[8] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[8] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[8] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[8], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[8], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[8], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[8], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[8] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[8] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[8] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[8] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[8], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[8], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[8], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[8], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[7] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[7] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[7] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[7] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$setup( posedge A2_0[7], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$setup( negedge A2_0[7], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$setup( posedge A2_0[7], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$setup( negedge A2_0[7], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[7] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[7] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[7] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[7] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$setup( posedge A2_0[7], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$setup( negedge A2_0[7], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$setup( posedge A2_0[7], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$setup( negedge A2_0[7], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[7] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[7] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[7] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[7] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[7], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[7], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[7], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[7], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[7] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[7] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[7] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[7] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[7], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[7], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[7], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[7], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[7] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[7] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[7] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[7] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[7], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[7], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[7], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[7], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[7] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[7] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[7] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[7] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[7], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[7], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[7], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[7], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[7] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[7] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[7] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[7] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[7], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[7], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[7], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[7], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[7] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[7] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[7] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[7] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[7], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[7], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[7], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[7], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[6] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[6] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[6] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[6] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$setup( posedge A2_0[6], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$setup( negedge A2_0[6], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$setup( posedge A2_0[6], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$setup( negedge A2_0[6], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[6] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[6] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[6] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[6] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$setup( posedge A2_0[6], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$setup( negedge A2_0[6], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$setup( posedge A2_0[6], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$setup( negedge A2_0[6], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[6] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[6] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[6] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[6] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[6], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[6], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[6], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[6], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[6] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[6] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[6] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[6] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[6], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[6], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[6], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[6], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[6] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[6] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[6] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[6] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[6], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[6], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[6], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[6], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[6] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[6] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[6] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[6] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[6], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[6], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[6], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[6], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[6] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[6] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[6] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[6] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[6], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[6], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[6], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[6], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[6] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[6] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[6] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[6] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[6], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[6], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[6], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[6], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[5] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[5] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[5] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[5] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$setup( posedge A2_0[5], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$setup( negedge A2_0[5], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$setup( posedge A2_0[5], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$setup( negedge A2_0[5], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[5] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[5] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[5] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[5] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$setup( posedge A2_0[5], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$setup( negedge A2_0[5], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$setup( posedge A2_0[5], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$setup( negedge A2_0[5], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[5] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[5] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[5] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[5] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[5], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[5], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[5], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[5], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[5] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[5] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[5] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[5] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[5], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[5], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[5], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[5], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[5] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[5] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[5] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[5] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[5], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[5], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[5], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[5], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[5] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[5] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[5] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[5] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[5], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[5], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[5], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[5], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[5] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[5] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[5] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[5] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[5], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[5], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[5], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[5], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[5] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[5] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[5] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[5] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[5], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[5], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[5], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[5], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[4] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[4] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[4] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[4] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$setup( posedge A2_0[4], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$setup( negedge A2_0[4], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$setup( posedge A2_0[4], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$setup( negedge A2_0[4], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[4] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[4] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[4] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[4] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$setup( posedge A2_0[4], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$setup( negedge A2_0[4], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$setup( posedge A2_0[4], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$setup( negedge A2_0[4], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[4] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[4] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[4] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[4] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[4], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[4], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[4], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[4], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[4] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[4] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[4] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[4] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[4], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[4], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[4], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[4], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[4] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[4] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[4] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[4] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[4], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[4], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[4], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[4], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[4] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[4] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[4] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[4] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[4], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[4], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[4], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[4], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[4] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[4] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[4] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[4] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[4], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[4], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[4], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[4], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[4] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[4] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[4] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[4] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[4], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[4], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[4], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[4], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[3] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[3] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[3] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[3] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$setup( posedge A2_0[3], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$setup( negedge A2_0[3], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$setup( posedge A2_0[3], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$setup( negedge A2_0[3], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[3] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[3] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[3] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[3] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$setup( posedge A2_0[3], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$setup( negedge A2_0[3], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$setup( posedge A2_0[3], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$setup( negedge A2_0[3], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[3] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[3] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[3] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[3] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[3], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[3], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[3], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[3], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[3] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[3] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[3] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[3] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[3], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[3], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[3], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[3], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[3] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[3] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[3] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[3] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[3], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[3], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[3], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[3], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[3] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[3] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[3] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[3] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[3], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[3], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[3], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[3], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[3] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[3] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[3] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[3] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[3], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[3], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[3], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[3], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[3] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[3] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[3] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[3] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[3], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[3], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[3], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[3], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[2] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[2] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[2] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[2] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$setup( posedge A2_0[2], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$setup( negedge A2_0[2], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$setup( posedge A2_0[2], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$setup( negedge A2_0[2], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[2] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[2] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[2] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[2] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$setup( posedge A2_0[2], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$setup( negedge A2_0[2], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$setup( posedge A2_0[2], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$setup( negedge A2_0[2], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[2] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[2] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[2] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[2] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[2], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[2], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[2], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[2], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[2] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[2] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[2] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[2] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[2], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[2], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[2], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[2], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[2] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[2] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[2] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[2] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[2], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[2], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[2], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[2], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[2] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[2] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[2] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[2] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[2], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[2], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[2], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[2], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[2] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[2] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[2] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[2] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[2], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[2], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[2], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[2], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[2] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[2] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[2] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[2] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[2], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[2], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[2], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[2], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[1] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[1] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[1] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[1] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$setup( posedge A2_0[1], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$setup( negedge A2_0[1], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$setup( posedge A2_0[1], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$setup( negedge A2_0[1], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[1] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[1] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[1] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[1] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$setup( posedge A2_0[1], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$setup( negedge A2_0[1], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$setup( posedge A2_0[1], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$setup( negedge A2_0[1], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[1] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[1] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[1] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[1] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[1], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[1], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[1], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[1], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[1] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[1] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[1] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[1] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[1], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[1], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[1], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[1], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[1] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[1] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[1] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[1] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[1], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[1], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[1], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[1], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[1] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[1] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[1] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[1] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[1], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[1], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[1], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[1], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[1] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[1] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[1] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[1] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[1], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[1], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[1], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[1], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[1] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[1] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[1] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[1] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[1], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[1], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[1], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[1], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[0] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[0] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[0] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[0] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$setup( posedge A2_0[0], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);
$setup( negedge A2_0[0], negedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_1, 0);


$setup( posedge A2_0[0], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);
$setup( negedge A2_0[0], posedge CLK2_1 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[0] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[0] &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[0] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[0] &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$setup( posedge A2_0[0], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);
$setup( negedge A2_0[0], negedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_1_0, 0);


$setup( posedge A2_0[0], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);
$setup( negedge A2_0[0], posedge CLK2_0 &&& ram01_addr2_18k_x36_hc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[0] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[0] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[0] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[0] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[0], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[0], negedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[0], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[0], posedge CLK2_1 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[0] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[0] &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[0] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[0] &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[0], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[0], negedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[0], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[0], posedge CLK2_0 &&& ram01_addr2_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge A2_0[0] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_0[0] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_0[0] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_0[0] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge A2_0[0], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge A2_0[0], negedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge A2_0[0], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge A2_0[0], posedge CLK2_1 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge A2_0[0] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[0] &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[0] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[0] &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge A2_0[0], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge A2_0[0], negedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge A2_0[0], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge A2_0[0], posedge CLK2_0 &&& ram01_addr2_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[0] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[0] &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[0] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[0] &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[0], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[0], negedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[0], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[0], posedge CLK2_0 &&& ram0_addr2_9k_x18_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge A2_0[0] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge A2_0[0] &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge A2_0[0] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge A2_0[0] &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$setup( posedge A2_0[0], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);
$setup( negedge A2_0[0], negedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_1_0, 0);


$setup( posedge A2_0[0], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);
$setup( negedge A2_0[0], posedge CLK2_0 &&& ram0_addr2_9k_x9_no_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[17] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[17] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[17] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[17] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[17], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[17], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[17], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[17], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[17], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[17], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[17], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[17], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[17], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[17], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[17], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[17], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[17] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[17], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[17], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[17], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[17], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[17] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[17] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[17] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[17] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[17], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[17], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[17], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[17], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[16] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[16] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[16] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[16] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[16], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[16], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[16], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[16], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[16], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[16], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[16], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[16], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[16], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[16], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[16], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[16], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[16] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[16], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[16], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[16], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[16], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[16] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[16] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[16] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[16] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[16], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[16], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[16], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[16], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[15] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[15] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[15] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[15] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[15], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[15], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[15], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[15], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[15], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[15], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[15], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[15], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[15], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[15], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[15], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[15], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[15] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[15], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[15], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[15], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[15], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[15] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[15] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[15] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[15] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[15], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[15], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[15], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[15], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[14] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[14] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[14] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[14] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[14], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[14], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[14], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[14], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[14], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[14], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[14], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[14], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[14], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[14], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[14], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[14], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[14] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[14], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[14], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[14], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[14], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[14] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[14] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[14] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[14] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[14], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[14], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[14], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[14], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[13] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[13] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[13] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[13] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[13], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[13], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[13], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[13], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[13], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[13], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[13], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[13], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[13], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[13], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[13], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[13], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[13] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[13], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[13], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[13], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[13], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[13] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[13] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[13] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[13] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[13], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[13], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[13], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[13], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[12] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[12] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[12] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[12] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[12], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[12], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[12], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[12], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[12], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[12], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[12], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[12], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[12], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[12], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[12], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[12], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[12] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[12], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[12], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[12], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[12], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[12] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[12] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[12] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[12] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[12], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[12], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[12], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[12], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[11] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[11] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[11] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[11] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[11], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[11], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[11], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[11], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[11], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[11], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[11], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[11], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[11], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[11], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[11], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[11], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[11] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[11], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[11], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[11], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[11], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[11] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[11] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[11] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[11] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[11], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[11], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[11], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[11], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[10] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[10] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[10] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[10] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[10], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[10], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[10], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[10], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[10], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[10], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[10], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[10], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[10], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[10], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[10], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[10], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[10] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[10], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[10], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[10], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[10], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[10] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[10] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[10] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[10] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[10], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[10], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[10], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[10], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[9] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[9] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[9] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[9] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[9], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[9], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[9], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[9], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[9], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[9], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[9], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[9], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[9], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[9], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[9], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[9], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[9] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[9], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[9], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[9], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[9], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[9] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[9] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[9] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[9] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[9], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[9], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[9], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[9], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[8] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[8] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[8] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[8] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[8], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[8], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[8], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[8], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[8], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[8], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[8], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[8], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[8], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[8], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[8], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[8], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[8], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[8], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[8], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[8], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[8], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[8], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[8], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[8], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[8] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[8], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[8], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[8], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[8], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[8] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[8] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[8] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[8] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[8], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[8], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[8], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[8], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[8] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[8] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[8] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[8] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[8], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[8], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[8], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[8], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[7] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[7] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[7] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[7] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[7], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[7], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[7], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[7], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[7], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[7], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[7], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[7], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[7], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[7], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[7], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[7], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[7], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[7], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[7], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[7], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[7], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[7], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[7], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[7], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[7] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[7], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[7], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[7], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[7], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[7] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[7] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[7] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[7] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[7], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[7], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[7], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[7], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[7] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[7] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[7] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[7] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[7], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[7], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[7], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[7], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[6] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[6] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[6] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[6] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[6], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[6], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[6], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[6], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[6], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[6], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[6], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[6], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[6], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[6], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[6], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[6], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[6], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[6], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[6], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[6], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[6], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[6], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[6], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[6], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[6] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[6], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[6], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[6], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[6], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[6] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[6] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[6] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[6] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[6], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[6], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[6], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[6], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[6] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[6] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[6] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[6] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[6], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[6], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[6], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[6], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[5] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[5] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[5] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[5] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[5], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[5], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[5], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[5], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[5], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[5], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[5], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[5], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[5], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[5], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[5], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[5], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[5], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[5], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[5], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[5], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[5], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[5], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[5], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[5], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[5] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[5], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[5], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[5], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[5], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[5] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[5] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[5] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[5] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[5], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[5], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[5], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[5], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[5] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[5] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[5] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[5] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[5], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[5], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[5], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[5], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[4] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[4] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[4] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[4] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[4], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[4], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[4], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[4], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[4], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[4], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[4], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[4], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[4], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[4], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[4], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[4], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[4], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[4], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[4], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[4], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[4], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[4], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[4], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[4], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[4] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[4], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[4], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[4], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[4], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[4] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[4] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[4] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[4] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[4], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[4], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[4], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[4], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[4] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[4] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[4] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[4] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[4], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[4], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[4], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[4], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[3] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[3] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[3] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[3] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[3], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[3], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[3], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[3], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[3], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[3], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[3], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[3], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[3], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[3], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[3], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[3], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[3], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[3], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[3], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[3], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[3], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[3], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[3], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[3], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[3] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[3], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[3], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[3], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[3], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[3] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[3] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[3] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[3] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[3], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[3], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[3], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[3], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[3] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[3] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[3] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[3] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[3], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[3], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[3], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[3], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[2] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[2] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[2] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[2] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[2], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[2], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[2], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[2], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[2], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[2], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[2], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[2], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[2], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[2], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[2], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[2], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[2], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[2], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[2], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[2], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[2], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[2], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[2], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[2], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[2] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[2], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[2], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[2], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[2], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[2] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[2] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[2] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[2] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[2], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[2], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[2], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[2], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[2] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[2] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[2] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[2] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[2], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[2], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[2], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[2], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[1] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[1] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[1] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[1] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[1], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[1], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[1], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[1], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[1], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[1], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[1], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[1], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[1], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[1], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[1], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[1], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[1], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[1], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[1], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[1], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[1], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[1], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[1], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[1], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[1] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[1], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[1], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[1], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[1], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[1] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[1] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[1] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[1] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[1], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[1], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[1], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[1], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[1] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[1] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[1] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[1] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[1], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[1], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[1], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[1], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[0] &&& fifo1_dir1_wd_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[0] &&& fifo1_dir1_wd_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[0] &&& fifo1_dir1_wd_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[0] &&& fifo1_dir1_wd_CLK2_0_1, 0);


$setup( posedge WD_1[0], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);
$setup( negedge WD_1[0], negedge CLK2_1 &&& fifo1_dir1_wd_CLK2_1_1, 0);


$setup( posedge WD_1[0], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);
$setup( negedge WD_1[0], posedge CLK2_1 &&& fifo1_dir1_wd_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$setup( posedge WD_1[0], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);
$setup( negedge WD_1[0], negedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_1_1, 0);


$setup( posedge WD_1[0], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);
$setup( negedge WD_1[0], posedge CLK1_1 &&& ram0_fifo_dir0_wd_18k_x36_hc_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[0], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[0], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[0], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[0], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[0], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[0], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[0], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[0], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x18_vc_con_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$setup( posedge WD_1[0], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);
$setup( negedge WD_1[0], negedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_1, 0);


$setup( posedge WD_1[0], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);
$setup( negedge WD_1[0], posedge CLK2_1 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WD_1[0] &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$setup( posedge WD_1[0], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);
$setup( negedge WD_1[0], negedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_1_0, 0);


$setup( posedge WD_1[0], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);
$setup( negedge WD_1[0], posedge CLK2_0 &&& ram0_fifo_dir0_wd_18k_x9_vc_con_CLK2_0_0, 0);


$hold( negedge CLK1_1, posedge WD_1[0] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[0] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[0] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[0] &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[0], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[0], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[0], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[0], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge WD_1[0] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WD_1[0] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WD_1[0] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WD_1[0] &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge WD_1[0], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge WD_1[0], negedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge WD_1[0], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge WD_1[0], posedge CLK1_1 &&& ram1_fifo_dir0_wd_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[9] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[9] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[9] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[9] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[9], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[9], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[9], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[9], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[8] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[8] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[8] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[8] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[8], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[8], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[8], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[8], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[8] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[8] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[8] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[8] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[8], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[8], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[8], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[8], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[7] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[7] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[7] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[7] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[7], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[7], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[7], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[7], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[7] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[7] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[7] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[7] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[7], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[7], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[7], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[7], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[6] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[6] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[6] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[6] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[6], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[6], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[6], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[6], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[6] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[6] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[6] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[6] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[6], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[6], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[6], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[6], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[5] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[5] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[5] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[5] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[5], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[5], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[5], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[5], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[5] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[5] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[5] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[5] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[5], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[5], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[5], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[5], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[4] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[4] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[4] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[4] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[4], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[4], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[4], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[4], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[4] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[4] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[4] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[4] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[4], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[4], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[4], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[4], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[3] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[3] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[3] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[3] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[3], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[3], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[3], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[3], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[3] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[3] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[3] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[3] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[3], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[3], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[3], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[3], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[2] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[2] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[2] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[2] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[2], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[2], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[2], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[2], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[2] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[2] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[2] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[2] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[2], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[2], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[2], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[2], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[1] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[1] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[1] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[1] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[1], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[1], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[1], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[1], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[1] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[1] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[1] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[1] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[1], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[1], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[1], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[1], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[0] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[0] &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[0] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[0] &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[0], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[0], negedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[0], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[0], posedge CLK1_1 &&& ram1_addr1_9k_x18_no_con_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge A1_1[0] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge A1_1[0] &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge A1_1[0] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge A1_1[0] &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$setup( posedge A1_1[0], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);
$setup( negedge A1_1[0], negedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_1_1, 0);


$setup( posedge A1_1[0], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);
$setup( negedge A1_1[0], posedge CLK1_1 &&& ram1_addr1_9k_x9_no_con_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);


$setup( posedge CS1_1, negedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);
$setup( negedge CS1_1, negedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);


$setup( posedge CS1_1, posedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);
$setup( negedge CS1_1, posedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);


$setup( posedge CS1_1, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);
$setup( negedge CS1_1, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);


$setup( posedge CS1_1, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);
$setup( negedge CS1_1, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);


$setup( posedge CS1_1, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);
$setup( negedge CS1_1, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);


$setup( posedge CS1_1, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);
$setup( negedge CS1_1, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);


$setup( posedge CS1_1, negedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);
$setup( negedge CS1_1, negedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);


$setup( posedge CS1_1, posedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);
$setup( negedge CS1_1, posedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_0_1, 0);


$setup( posedge CS1_1, negedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_1_1, 0);
$setup( negedge CS1_1, negedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_1_1, 0);


$setup( posedge CS1_1, posedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_0_1, 0);
$setup( negedge CS1_1, posedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_0_1, 0);


$setup( posedge CS1_1, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_1_1, 0);
$setup( negedge CS1_1, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_1_1, 0);


$setup( posedge CS1_1, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_0_1, 0);
$setup( negedge CS1_1, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_0_1, 0);


$setup( posedge CS1_1, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_1_1, 0);
$setup( negedge CS1_1, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_1_1, 0);


$setup( posedge CS1_1, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_0_1, 0);
$setup( negedge CS1_1, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_0_1, 0);


$setup( posedge CS1_1, negedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_1_1, 0);
$setup( negedge CS1_1, negedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_1_1, 0);


$setup( posedge CS1_1, posedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_0_1, 0);
$setup( negedge CS1_1, posedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge WEN1_1[1] &&& ram1_wen_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WEN1_1[1] &&& ram1_wen_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WEN1_1[1] &&& ram1_wen_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WEN1_1[1] &&& ram1_wen_CLK2_0_1, 0);


$setup( posedge WEN1_1[1], negedge CLK2_1 &&& ram1_wen_CLK2_1_1, 0);
$setup( negedge WEN1_1[1], negedge CLK2_1 &&& ram1_wen_CLK2_1_1, 0);


$setup( posedge WEN1_1[1], posedge CLK2_1 &&& ram1_wen_CLK2_0_1, 0);
$setup( negedge WEN1_1[1], posedge CLK2_1 &&& ram1_wen_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WEN1_1[1] &&& ram1_wen_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WEN1_1[1] &&& ram1_wen_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WEN1_1[1] &&& ram1_wen_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WEN1_1[1] &&& ram1_wen_CLK1_0_1, 0);


$setup( posedge WEN1_1[1], negedge CLK1_1 &&& ram1_wen_CLK1_1_1, 0);
$setup( negedge WEN1_1[1], negedge CLK1_1 &&& ram1_wen_CLK1_1_1, 0);


$setup( posedge WEN1_1[1], posedge CLK1_1 &&& ram1_wen_CLK1_0_1, 0);
$setup( negedge WEN1_1[1], posedge CLK1_1 &&& ram1_wen_CLK1_0_1, 0);


$hold( negedge CLK2_0, posedge WEN1_1[1] &&& ram1_wen_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WEN1_1[1] &&& ram1_wen_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WEN1_1[1] &&& ram1_wen_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WEN1_1[1] &&& ram1_wen_CLK2_0_0, 0);


$setup( posedge WEN1_1[1], negedge CLK2_0 &&& ram1_wen_CLK2_1_0, 0);
$setup( negedge WEN1_1[1], negedge CLK2_0 &&& ram1_wen_CLK2_1_0, 0);


$setup( posedge WEN1_1[1], posedge CLK2_0 &&& ram1_wen_CLK2_0_0, 0);
$setup( negedge WEN1_1[1], posedge CLK2_0 &&& ram1_wen_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge WEN1_1[0] &&& ram1_wen_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge WEN1_1[0] &&& ram1_wen_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge WEN1_1[0] &&& ram1_wen_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge WEN1_1[0] &&& ram1_wen_CLK2_0_1, 0);


$setup( posedge WEN1_1[0], negedge CLK2_1 &&& ram1_wen_CLK2_1_1, 0);
$setup( negedge WEN1_1[0], negedge CLK2_1 &&& ram1_wen_CLK2_1_1, 0);


$setup( posedge WEN1_1[0], posedge CLK2_1 &&& ram1_wen_CLK2_0_1, 0);
$setup( negedge WEN1_1[0], posedge CLK2_1 &&& ram1_wen_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge WEN1_1[0] &&& ram1_wen_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge WEN1_1[0] &&& ram1_wen_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge WEN1_1[0] &&& ram1_wen_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge WEN1_1[0] &&& ram1_wen_CLK1_0_1, 0);


$setup( posedge WEN1_1[0], negedge CLK1_1 &&& ram1_wen_CLK1_1_1, 0);
$setup( negedge WEN1_1[0], negedge CLK1_1 &&& ram1_wen_CLK1_1_1, 0);


$setup( posedge WEN1_1[0], posedge CLK1_1 &&& ram1_wen_CLK1_0_1, 0);
$setup( negedge WEN1_1[0], posedge CLK1_1 &&& ram1_wen_CLK1_0_1, 0);


$hold( negedge CLK2_0, posedge WEN1_1[0] &&& ram1_wen_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge WEN1_1[0] &&& ram1_wen_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge WEN1_1[0] &&& ram1_wen_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge WEN1_1[0] &&& ram1_wen_CLK2_0_0, 0);


$setup( posedge WEN1_1[0], negedge CLK2_0 &&& ram1_wen_CLK2_1_0, 0);
$setup( negedge WEN1_1[0], negedge CLK2_0 &&& ram1_wen_CLK2_1_0, 0);


$setup( posedge WEN1_1[0], posedge CLK2_0 &&& ram1_wen_CLK2_0_0, 0);
$setup( negedge WEN1_1[0], posedge CLK2_0 &&& ram1_wen_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);


$setup( posedge CS2_1, negedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);
$setup( negedge CS2_1, negedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);


$setup( posedge CS2_1, posedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);
$setup( negedge CS2_1, posedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);


$setup( posedge CS2_1, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);
$setup( negedge CS2_1, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);


$setup( posedge CS2_1, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);
$setup( negedge CS2_1, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);


$setup( posedge CS2_1, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);
$setup( negedge CS2_1, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_1_1, 0);


$setup( posedge CS2_1, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);
$setup( negedge CS2_1, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);


$setup( posedge CS2_1, negedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);
$setup( negedge CS2_1, negedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_1_1, 0);


$setup( posedge CS2_1, posedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);
$setup( negedge CS2_1, posedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat1_hc_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_0_1, 0);


$setup( posedge CS2_1, negedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_1_1, 0);
$setup( negedge CS2_1, negedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_1_1, 0);


$setup( posedge CS2_1, posedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_0_1, 0);
$setup( negedge CS2_1, posedge CLK2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS2_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_0_1, 0);


$setup( posedge CS2_1, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_1_1, 0);
$setup( negedge CS2_1, negedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_1_1, 0);


$setup( posedge CS2_1, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_0_1, 0);
$setup( negedge CS2_1, posedge CLK1_1 &&& fifo0_dir1_cs1_cs2_ram1_concat0_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_0_1, 0);


$setup( posedge CS2_1, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_1_1, 0);
$setup( negedge CS2_1, negedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_1_1, 0);


$setup( posedge CS2_1, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_0_1, 0);
$setup( negedge CS2_1, posedge CLK2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge CS2_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_0_1, 0);


$setup( posedge CS2_1, negedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_1_1, 0);
$setup( negedge CS2_1, negedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_1_1, 0);


$setup( posedge CS2_1, posedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_0_1, 0);
$setup( negedge CS2_1, posedge CLK1_1 &&& fifo0_dir0_cs1_cs2_ram1_concat0_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[9] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[9] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[9] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[9] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[9], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[9], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[9], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[9], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[8] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[8] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[8] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[8] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[8], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[8], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[8], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[8], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[8] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[8] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[8] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[8] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[8], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[8], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[8], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[8], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[7] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[7] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[7] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[7] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[7], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[7], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[7], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[7], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[7] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[7] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[7] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[7] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[7], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[7], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[7], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[7], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[6] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[6] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[6] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[6] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[6], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[6], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[6], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[6], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[6] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[6] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[6] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[6] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[6], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[6], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[6], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[6], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[5] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[5] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[5] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[5] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[5], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[5], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[5], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[5], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[5] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[5] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[5] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[5] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[5], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[5], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[5], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[5], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[4] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[4] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[4] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[4] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[4], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[4], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[4], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[4], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[4] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[4] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[4] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[4] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[4], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[4], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[4], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[4], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[3] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[3] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[3] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[3] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[3], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[3], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[3], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[3], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[3] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[3] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[3] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[3] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[3], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[3], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[3], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[3], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[2] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[2] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[2] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[2] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[2], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[2], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[2], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[2], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[2] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[2] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[2] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[2] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[2], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[2], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[2], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[2], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[1] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[1] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[1] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[1] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[1], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[1], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[1], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[1], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[1] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[1] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[1] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[1] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[1], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[1], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[1], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[1], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[0] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[0] &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[0] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[0] &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[0], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[0], negedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[0], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[0], posedge CLK2_1 &&& ram1_addr2_9k_x18_no_con_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge A2_1[0] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge A2_1[0] &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge A2_1[0] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge A2_1[0] &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$setup( posedge A2_1[0], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);
$setup( negedge A2_1[0], negedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_1_1, 0);


$setup( posedge A2_1[0], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);
$setup( negedge A2_1[0], posedge CLK2_1 &&& ram1_add2r_9k_x9_no_con_CLK2_0_1, 0);


$hold( negedge CLK1_1, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_1, 0);


$setup( posedge P1_0, negedge CLK1_1 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_1, 0);
$setup( negedge P1_0, negedge CLK1_1 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_1, 0);


$setup( posedge P1_0, posedge CLK1_1 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_1, 0);
$setup( negedge P1_0, posedge CLK1_1 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_0, 0);


$setup( posedge P1_0, negedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_0, 0);
$setup( negedge P1_0, negedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_1_0, 0);


$setup( posedge P1_0, posedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_0, 0);
$setup( negedge P1_0, posedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_1, 0);


$setup( posedge P1_0, negedge CLK1_1 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_1, 0);
$setup( negedge P1_0, negedge CLK1_1 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_1, 0);


$setup( posedge P1_0, posedge CLK1_1 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_1, 0);
$setup( negedge P1_0, posedge CLK1_1 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_0, 0);


$setup( posedge P1_0, negedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_0, 0);
$setup( negedge P1_0, negedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_1_0, 0);


$setup( posedge P1_0, posedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_0, 0);
$setup( negedge P1_0, posedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_1, 0);


$setup( posedge P1_0, negedge CLK1_1 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_1, 0);
$setup( negedge P1_0, negedge CLK1_1 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_1, 0);


$setup( posedge P1_0, posedge CLK1_1 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_1, 0);
$setup( negedge P1_0, posedge CLK1_1 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_0, 0);


$setup( posedge P1_0, negedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_0, 0);
$setup( negedge P1_0, negedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_1_0, 0);


$setup( posedge P1_0, posedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_0, 0);
$setup( negedge P1_0, posedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_1, 0);


$setup( posedge P1_0, negedge CLK1_1 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_1, 0);
$setup( negedge P1_0, negedge CLK1_1 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_1, 0);


$setup( posedge P1_0, posedge CLK1_1 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_1, 0);
$setup( negedge P1_0, posedge CLK1_1 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_1, 0);


$hold( negedge CLK1_0, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_0, 0);


$setup( posedge P1_0, negedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_0, 0);
$setup( negedge P1_0, negedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_1_0, 0);


$setup( posedge P1_0, posedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_0, 0);
$setup( negedge P1_0, posedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge P1_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK1_0_0, 0);


$setup( posedge P1_0, negedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK1_1_0, 0);
$setup( negedge P1_0, negedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK1_1_0, 0);


$setup( posedge P1_0, posedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK1_0_0, 0);
$setup( negedge P1_0, posedge CLK1_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK1_0_0, 0);


$hold( negedge CLK1_0, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK1_1_0, 0);
$hold( negedge CLK1_0, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK1_1_0, 0);


$hold( posedge CLK1_0, posedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK1_0_0, 0);
$hold( posedge CLK1_0, negedge P1_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK1_0_0, 0);


$setup( posedge P1_0, negedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK1_1_0, 0);
$setup( negedge P1_0, negedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK1_1_0, 0);


$setup( posedge P1_0, posedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK1_0_0, 0);
$setup( negedge P1_0, posedge CLK1_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK1_0_0, 0);


$hold( negedge CLK1_1, posedge P1_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge P1_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge P1_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge P1_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_0_1, 0);


$setup( posedge P1_1, negedge CLK1_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_1_1, 0);
$setup( negedge P1_1, negedge CLK1_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_1_1, 0);


$setup( posedge P1_1, posedge CLK1_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_0_1, 0);
$setup( negedge P1_1, posedge CLK1_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge P1_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge P1_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge P1_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge P1_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_0_1, 0);


$setup( posedge P1_1, negedge CLK1_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_1_1, 0);
$setup( negedge P1_1, negedge CLK1_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_1_1, 0);


$setup( posedge P1_1, posedge CLK1_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_0_1, 0);
$setup( negedge P1_1, posedge CLK1_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge P1_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge P1_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge P1_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge P1_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK1_0_1, 0);


$setup( posedge P1_1, negedge CLK1_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK1_1_1, 0);
$setup( negedge P1_1, negedge CLK1_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK1_1_1, 0);


$setup( posedge P1_1, posedge CLK1_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK1_0_1, 0);
$setup( negedge P1_1, posedge CLK1_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK1_0_1, 0);


$hold( negedge CLK1_1, posedge P1_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK1_1_1, 0);
$hold( negedge CLK1_1, negedge P1_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK1_1_1, 0);


$hold( posedge CLK1_1, posedge P1_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK1_0_1, 0);
$hold( posedge CLK1_1, negedge P1_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK1_0_1, 0);


$setup( posedge P1_1, negedge CLK1_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK1_1_1, 0);
$setup( negedge P1_1, negedge CLK1_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK1_1_1, 0);


$setup( posedge P1_1, posedge CLK1_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK1_0_1, 0);
$setup( negedge P1_1, posedge CLK1_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK1_0_1, 0);


$hold( negedge CLK2_1, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_1, 0);


$setup( posedge P2_0, negedge CLK2_1 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_1, 0);
$setup( negedge P2_0, negedge CLK2_1 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_1, 0);


$setup( posedge P2_0, posedge CLK2_1 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_1, 0);
$setup( negedge P2_0, posedge CLK2_1 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_0, 0);


$setup( posedge P2_0, negedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_0, 0);
$setup( negedge P2_0, negedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_1_0, 0);


$setup( posedge P2_0, posedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_0, 0);
$setup( negedge P2_0, posedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_hc_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_1, 0);


$setup( posedge P2_0, negedge CLK2_1 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_1, 0);
$setup( negedge P2_0, negedge CLK2_1 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_1, 0);


$setup( posedge P2_0, posedge CLK2_1 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_1, 0);
$setup( negedge P2_0, posedge CLK2_1 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_0, 0);


$setup( posedge P2_0, negedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_0, 0);
$setup( negedge P2_0, negedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_1_0, 0);


$setup( posedge P2_0, posedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_0, 0);
$setup( negedge P2_0, posedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_hc_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_1, 0);


$setup( posedge P2_0, negedge CLK2_1 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_1, 0);
$setup( negedge P2_0, negedge CLK2_1 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_1, 0);


$setup( posedge P2_0, posedge CLK2_1 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_1, 0);
$setup( negedge P2_0, posedge CLK2_1 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_0, 0);


$setup( posedge P2_0, negedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_0, 0);
$setup( negedge P2_0, negedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_1_0, 0);


$setup( posedge P2_0, posedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_0, 0);
$setup( negedge P2_0, posedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat1_vc_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_1, 0);


$setup( posedge P2_0, negedge CLK2_1 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_1, 0);
$setup( negedge P2_0, negedge CLK2_1 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_1, 0);


$setup( posedge P2_0, posedge CLK2_1 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_1, 0);
$setup( negedge P2_0, posedge CLK2_1 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_1, 0);


$hold( negedge CLK2_0, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_0, 0);


$setup( posedge P2_0, negedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_0, 0);
$setup( negedge P2_0, negedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_1_0, 0);


$setup( posedge P2_0, posedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_0, 0);
$setup( negedge P2_0, posedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat1_vc_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge P2_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK2_0_0, 0);


$setup( posedge P2_0, negedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK2_1_0, 0);
$setup( negedge P2_0, negedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK2_1_0, 0);


$setup( posedge P2_0, posedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK2_0_0, 0);
$setup( negedge P2_0, posedge CLK2_0 &&& fifo0_dir1_p1_p2_ram0_concat0_CLK2_0_0, 0);


$hold( negedge CLK2_0, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK2_1_0, 0);
$hold( negedge CLK2_0, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK2_1_0, 0);


$hold( posedge CLK2_0, posedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK2_0_0, 0);
$hold( posedge CLK2_0, negedge P2_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK2_0_0, 0);


$setup( posedge P2_0, negedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK2_1_0, 0);
$setup( negedge P2_0, negedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK2_1_0, 0);


$setup( posedge P2_0, posedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK2_0_0, 0);
$setup( negedge P2_0, posedge CLK2_0 &&& fifo0_dir0_p1_p2_ram0_concat0_CLK2_0_0, 0);


$hold( negedge CLK2_1, posedge P2_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge P2_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge P2_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge P2_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_0_1, 0);


$setup( posedge P2_1, negedge CLK2_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_1_1, 0);
$setup( negedge P2_1, negedge CLK2_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_1_1, 0);


$setup( posedge P2_1, posedge CLK2_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_0_1, 0);
$setup( negedge P2_1, posedge CLK2_1 &&& fifo0_dir1_p1_p2_ram1_concat1_hc_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge P2_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge P2_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge P2_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge P2_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_0_1, 0);


$setup( posedge P2_1, negedge CLK2_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_1_1, 0);
$setup( negedge P2_1, negedge CLK2_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_1_1, 0);


$setup( posedge P2_1, posedge CLK2_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_0_1, 0);
$setup( negedge P2_1, posedge CLK2_1 &&& fifo0_dir0_p1_p2_ram1_concat1_hc_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge P2_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge P2_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge P2_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge P2_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK2_0_1, 0);


$setup( posedge P2_1, negedge CLK2_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK2_1_1, 0);
$setup( negedge P2_1, negedge CLK2_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK2_1_1, 0);


$setup( posedge P2_1, posedge CLK2_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK2_0_1, 0);
$setup( negedge P2_1, posedge CLK2_1 &&& fifo0_dir1_p1_p2_ram1_concat0_CLK2_0_1, 0);


$hold( negedge CLK2_1, posedge P2_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK2_1_1, 0);
$hold( negedge CLK2_1, negedge P2_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK2_1_1, 0);


$hold( posedge CLK2_1, posedge P2_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK2_0_1, 0);
$hold( posedge CLK2_1, negedge P2_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK2_0_1, 0);


$setup( posedge P2_1, negedge CLK2_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK2_1_1, 0);
$setup( negedge P2_1, negedge CLK2_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK2_1_1, 0);


$setup( posedge P2_1, posedge CLK2_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK2_0_1, 0);
$setup( negedge P2_1, posedge CLK2_1 &&& fifo0_dir0_p1_p2_ram1_concat0_CLK2_0_1, 0);


$recovery( posedge CLK1_0, negedge CLK2_0 &&& fifo0_dir1_sync_CLK2_1_0, 0);
$recovery( negedge CLK1_0, negedge CLK2_0 &&& fifo0_dir1_sync_CLK2_1_0, 0);


$recovery( posedge CLK1_0, posedge CLK2_0 &&& fifo0_dir1_sync_CLK2_0_0, 0);
$recovery( negedge CLK1_0, posedge CLK2_0 &&& fifo0_dir1_sync_CLK2_0_0, 0);


$recovery( posedge CLK1_0, negedge CLK2_0 &&& fifo0_dir0_sync_CLK2_1_0, 0);
$recovery( negedge CLK1_0, negedge CLK2_0 &&& fifo0_dir0_sync_CLK2_1_0, 0);


$recovery( posedge CLK1_0, posedge CLK2_0 &&& fifo0_dir0_sync_CLK2_0_0, 0);
$recovery( negedge CLK1_0, posedge CLK2_0 &&& fifo0_dir0_sync_CLK2_0_0, 0);


$recovery( posedge CLK1_1, negedge CLK2_1 &&& fifo1_dir1_sync_CLK2_1_1, 0);
$recovery( negedge CLK1_1, negedge CLK2_1 &&& fifo1_dir1_sync_CLK2_1_1, 0);


$recovery( posedge CLK1_1, posedge CLK2_1 &&& fifo1_dir1_sync_CLK2_0_1, 0);
$recovery( negedge CLK1_1, posedge CLK2_1 &&& fifo1_dir1_sync_CLK2_0_1, 0);


$recovery( posedge CLK1_1, negedge CLK2_1 &&& fifo1_dir0_sync_CLK2_1_1, 0);
$recovery( negedge CLK1_1, negedge CLK2_1 &&& fifo1_dir0_sync_CLK2_1_1, 0);


$recovery( posedge CLK1_1, posedge CLK2_1 &&& fifo1_dir0_sync_CLK2_0_1, 0);
$recovery( negedge CLK1_1, posedge CLK2_1 &&& fifo1_dir0_sync_CLK2_0_1, 0);


$recovery( posedge CLK2_0, negedge CLK1_0 &&& fifo0_dir1_sync_CLK1_1_0, 0);
$recovery( negedge CLK2_0, negedge CLK1_0 &&& fifo0_dir1_sync_CLK1_1_0, 0);


$recovery( posedge CLK2_0, posedge CLK1_0 &&& fifo0_dir1_sync_CLK1_0_0, 0);
$recovery( negedge CLK2_0, posedge CLK1_0 &&& fifo0_dir1_sync_CLK1_0_0, 0);


$recovery( posedge CLK2_0, negedge CLK1_0 &&& fifo0_dir0_sync_CLK1_1_0, 0);
$recovery( negedge CLK2_0, negedge CLK1_0 &&& fifo0_dir0_sync_CLK1_1_0, 0);


$recovery( posedge CLK2_0, posedge CLK1_0 &&& fifo0_dir0_sync_CLK1_0_0, 0);
$recovery( negedge CLK2_0, posedge CLK1_0 &&& fifo0_dir0_sync_CLK1_0_0, 0);


$recovery( posedge CLK2_1, negedge CLK1_1 &&& fifo1_dir1_sync_CLK1_1_1, 0);
$recovery( negedge CLK2_1, negedge CLK1_1 &&& fifo1_dir1_sync_CLK1_1_1, 0);


$recovery( posedge CLK2_1, posedge CLK1_1 &&& fifo1_dir1_sync_CLK1_0_1, 0);
$recovery( negedge CLK2_1, posedge CLK1_1 &&& fifo1_dir1_sync_CLK1_0_1, 0);


$recovery( posedge CLK2_1, negedge CLK1_1 &&& fifo1_dir0_sync_CLK1_1_1, 0);
$recovery( negedge CLK2_1, negedge CLK1_1 &&& fifo1_dir0_sync_CLK1_1_1, 0);


$recovery( posedge CLK2_1, posedge CLK1_1 &&& fifo1_dir0_sync_CLK1_0_1, 0);
$recovery( negedge CLK2_1, posedge CLK1_1 &&& fifo1_dir0_sync_CLK1_0_1, 0);


endspecify
/*********************************/

//pragma synthesis_on
endmodule

//--------------------RAM8K...........................

// P_MUX3 cell -----------------------------------------------------------------

module P_MUX3( A, B, C, D, S, T, E, Z );
input A, B, C, D, S, E, T;
output Z;

udpmux3 QL2 ( Z, A, B, C, D, E, S, T );

specify
   (A => Z) = 0;
   (B => Z) = 0;
   (C => Z) = 0;
   (D => Z) = 0;
   (E => Z) = 0;
   (S => Z) = 0;
   (T => Z) = 0;
endspecify

endmodule

primitive udpmux3(Z, A, B, C, D, E, S, T);
   output Z;
   input A, B, C, D, E, S, T;
   table
   // A  B  C  D  E     S  T   :    Z
      1  ?  ?  ?  ?     0  0   :    1  ;
      0  ?  ?  ?  ?     0  0   :    0  ;
      ?  0  ?  ?  ?     0  1   :    0  ;
      ?  1  ?  ?  ?     0  1   :    1  ;
      ?  ?  0  ?  ?     1  0   :    0  ;
      ?  ?  1  ?  ?     1  0   :    1  ;
      ?  ?  ?  0  ?     1  1   :    0  ;
      ?  ?  ?  1  ?     1  1   :    1  ;
   endtable
endprimitive // udpmux3

// P_MUX2 cell -----------------------------------------------------------------


module P_MUX2( A, B, C, D, S, Z);
input A, B, C, D, S;
output Z;

udpmux2 QL1 ( Z, A, B, C, D, S );

specify
   (A => Z) = 0;
   (B => Z) = 0;
   (C => Z) = 0;
   (D => Z) = 0;
   (S => Z) = 0;
endspecify

endmodule // P_MUX2

// P_BUF cell -----------------------------------------------------------------

module P_BUF( A, Z);
input A;
output Z;

buf QL1 (Z, A);

specify
   (A => Z) = 0;
endspecify

endmodule

primitive udpmux2(Z, A, B, C, D, S);
   output Z;
   input A, B, C, D, S;
   table
      // A  B  C  D  S   :    Z
         1  0  ?  ?  0   :    1  ;
         0  ?  ?  ?  0   :    0  ;
         ?  1  ?  ?  0   :    0  ;
         ?  ?  1  0  1   :    1  ;
         ?  ?  0  ?  1   :    0  ;
         ?  ?  ?  1  1   :    0  ;
// Reduce pessimism
         1  0  1  0  ?   :    1  ;
         0  ?  0  ?  ?   :    0  ;
         0  ?  ?  1  ?   :    0  ; // new
         ?  1  ?  1  ?   :    0  ;
         ?  1  0  ?  ?   :    0  ; // new
   endtable
endprimitive // udpmux2

primitive udpand6(Z, A, B, C, D, E, F);
   output Z;
   input A, B, C, D, E, F;
   table
      // A  B  C  D  E  F  :  Z
         1  0  1  0  1  0  :  1  ;
         0  ?  ?  ?  ?  ?  :  0  ;
         ?  1  ?  ?  ?  ?  :  0  ;
         ?  ?  0  ?  ?  ?  :  0  ;
         ?  ?  ?  1  ?  ?  :  0  ;
         ?  ?  ?  ?  0  ?  :  0  ;
         ?  ?  ?  ?  ?  1  :  0  ;
   endtable
endprimitive // udpand6

module P_AND6( A, B, C, D, E, F, Z );
input A, B, C, D, E, F;
output Z;

udpand6 QL1 ( Z, A, B, C, D, E, F );

specify
   (A => Z) = 0;
   (B => Z) = 0;
   (C => Z) = 0;
   (D => Z) = 0;
   (E => Z) = 0;
   (F => Z) = 0;
endspecify

endmodule // P_AND6

module P_MULT(
		input [31:0] Amult,
		input [31:0] Bmult,
		output [63:0] Cmult,
		input [1:0] Valid_mult,
		input sel_mul_32x32
);

wire [31:0] Amult_int;
wire [31:0] Bmult_int;
wire [1:0] Valid_mult_int;	
wire sel_mul_32x32_int;

buf Amult_buf[31:0] (Amult_int,Amult);
buf Bmult_buf[31:0] (Bmult_int,Bmult);
buf Valid_mult_buf[1:0] (Valid_mult_int,Valid_mult);	
buf sel_mul_32x32_buf (sel_mul_32x32_int,sel_mul_32x32);

qlal4s3_mult_cell_macro inst_qlal4s3_mult_cell (
		 .Amult(Amult_int),
		 .Bmult(Bmult_int),
		 .Valid_mult(Valid_mult_int),
		 .sel_mul_32x32(sel_mul_32x32_int),
		 .Cmult(Cmult)
		);

specify

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[0]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[0]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[0]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[0]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[1]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[1]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[1]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[1]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[1]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[1]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[1]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[1]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[2]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[3]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[4]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[5]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[6]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[7]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[8]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[9]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[10]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[11]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[12]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[13]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[14]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[15]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[16]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[17]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[18]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[19]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[20]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[21]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[22]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[23]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[24]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[25]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[26]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[27]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[28]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[29]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[30]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[15] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[14] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[13] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[12] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[11] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[10] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[9] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[8] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[7] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[6] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[5] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[4] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[3] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[2] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[1] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[0] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[15] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[14] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[13] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[12] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[11] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[10] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[9] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[8] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[7] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[6] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[5] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[4] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[3] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[2] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[1] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[0] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[31]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[32]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[32]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[32]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[33]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[33]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[33]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[33]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[33]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[34]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[34]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[34]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[34]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[34]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[34]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[34]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[35]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[35]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[35]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[35]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[35]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[35]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[35]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[35]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[35]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[36]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[36]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[37]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[37]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[38]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[38]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[39]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[39]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[40]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[40]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[41]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[41]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[42]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[42]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[43]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[43]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[44]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[44]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[45]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[45]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[46]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[46]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[47]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[47]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[48]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[48]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[49]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[49]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[50]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[50]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[51]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[51]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[52]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[52]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[53]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[53]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[54]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[54]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[55]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[55]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[56]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[56]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[57]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[57]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[58]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[58]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[59]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[59]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[60]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[60]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[61]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[61]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[62]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[62]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[31] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[31] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[30] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[30] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[29] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[29] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[28] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[28] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[27] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[27] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[26] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[26] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[25] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[25] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[24] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[24] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[23] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[23] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[22] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[22] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[21] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[21] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[20] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[20] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[19] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[19] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[18] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[18] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[17] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[17] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Bmult[16] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[16] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[15] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[14] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[13] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[12] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[11] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[10] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[9] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[8] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[7] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[6] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[5] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[4] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[3] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[2] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[1] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Bmult[0] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[31] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[31] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[30] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[30] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[29] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[29] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[28] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[28] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[27] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[27] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[26] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[26] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[25] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[25] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[24] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[24] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[23] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[23] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[22] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[22] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[21] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[21] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[20] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[20] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[19] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[19] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[18] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[18] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[17] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[17] => Cmult[63]) = (0,0);

if (Valid_mult[1] == 1'b1  && sel_mul_32x32 == 1'b0)
(Amult[16] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[16] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[15] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[14] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[13] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[12] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[11] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[10] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[9] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[8] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[7] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[6] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[5] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[4] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[3] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[2] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[1] => Cmult[63]) = (0,0);

if (Valid_mult[0] == 1'b1  && sel_mul_32x32 == 1'b1)
(Amult[0] => Cmult[63]) = (0,0);

endspecify

endmodule /* qlal4s3_mult_cell*/

module P_ASSPTMRB(
					WB_CLK, WBs_ACK, WBs_RD_DAT, WBs_BYTE_STB, WBs_CYC, WBs_WE,
					WBs_RD, WBs_STB, WBs_ADR, SDMA_Req, SDMA_Sreq, SDMA_Done,
					SDMA_Active, FB_msg_out, FB_Int_Clr, FB_Start, FB_Busy,
					WB_RST, Sys_PKfb_Rst, Sys_Clk0, Sys_Clk0_Rst, Sys_Clk1,
					Sys_Clk1_Rst, Sys_Pclk, Sys_Pclk_Rst, Sys_PKfb_Clk, 
					FB_PKfbData, WBs_WR_DAT, FB_PKfbPush, FB_PKfbSOF, FB_PKfbEOF,
					Sensor_Int, FB_PKfbOverflow, TimeStamp, Sys_PSel, SPIm_Paddr,
					SPIm_PEnable, SPIm_PWrite, SPIm_PWdata, SPIm_PReady, 
					SPIm_PSlvErr, SPIm_Prdata, Device_ID, FBIO_In_En, FBIO_Out,
					FBIO_Out_En, FBIO_In, Device_ID_6S, Device_ID_4S, SPIm_PWdata_26S, 
					SPIm_PWdata_24S, SPIm_PWdata_14S, SPIm_PWdata_11S, SPIm_PWdata_0S, 
					SPIm_Paddr_8S, SPIm_Paddr_6S, FB_PKfbPush_1S, FB_PKfbData_31S, 
					FB_PKfbData_21S, FB_PKfbData_19S, FB_PKfbData_9S, FB_PKfbData_6S,
					Sys_PKfb_ClkS, FB_BusyS, WB_CLKS, SFBIO);
			
input	WB_CLK;
input	WBs_ACK;
input	[31:0]WBs_RD_DAT;
output	[3:0]WBs_BYTE_STB;
output	WBs_CYC;
output	WBs_WE;
output	WBs_RD;
output	WBs_STB;
output	[16:0]WBs_ADR;
input	[3:0]SDMA_Req;
input	[3:0]SDMA_Sreq;
output	[3:0]SDMA_Done;
output	[3:0]SDMA_Active;
input	[3:0]FB_msg_out;
input	[7:0]FB_Int_Clr;
output	FB_Start;
input	FB_Busy;
output	WB_RST;
output	Sys_PKfb_Rst;
output	Sys_Clk0;
output	Sys_Clk0_Rst;
output	Sys_Clk1;
output	Sys_Clk1_Rst;
output	Sys_Pclk;
output	Sys_Pclk_Rst;
input	Sys_PKfb_Clk;
input	[31:0]FB_PKfbData;
output	[31:0]WBs_WR_DAT;
input	[3:0]FB_PKfbPush;
input	FB_PKfbSOF;
input	FB_PKfbEOF;
output	[7:0]Sensor_Int;
output	FB_PKfbOverflow;
output	[23:0]TimeStamp;
input	Sys_PSel;
input	[15:0]SPIm_Paddr;
input	SPIm_PEnable;
input	SPIm_PWrite;
input	[31:0]SPIm_PWdata;
output	SPIm_PReady;
output	SPIm_PSlvErr;
output	[31:0]SPIm_Prdata;
input	[15:0]Device_ID;
input	[13:0]FBIO_In_En;
input	[13:0]FBIO_Out;
input	[13:0]FBIO_Out_En;
output	[13:0]FBIO_In;
inout 	[13:0]SFBIO;

input   Device_ID_6S; 
input   Device_ID_4S; 
input   SPIm_PWdata_26S; 
input   SPIm_PWdata_24S;  
input   SPIm_PWdata_14S; 
input   SPIm_PWdata_11S; 
input   SPIm_PWdata_0S; 
input   SPIm_Paddr_8S; 
input   SPIm_Paddr_6S; 
input   FB_PKfbPush_1S; 
input   FB_PKfbData_31S; 
input   FB_PKfbData_21S;
input   FB_PKfbData_19S;
input   FB_PKfbData_9S;
input   FB_PKfbData_6S;
input   Sys_PKfb_ClkS;
input   FB_BusyS;
input	WB_CLKS;

wire	WB_CLK_int;
wire	WBs_ACK_int;
wire	[31:0]WBs_RD_DAT_int;
wire	[3:0]SDMA_Req_int;
wire	[3:0]SDMA_Sreq_int;
wire	[3:0]FB_msg_out_int;
wire	[7:0]FB_Int_Clr_int;
wire	FB_Busy_int;
wire	Sys_PKfb_Clk_int;
wire	[31:0]FB_PKfbData_int;
wire	[3:0]FB_PKfbPush_int;
wire	FB_PKfbSOF_int;
wire	FB_PKfbEOF_int;
wire	Sys_PSel_int;
wire	[15:0]SPIm_Paddr_int;
wire	SPIm_PEnable_int;
wire	SPIm_PWrite_int;
wire	[31:0]SPIm_PWdata_int;
wire	[15:0]Device_ID_int;
wire	[13:0]FBIO_In_En_int;
wire	[13:0]FBIO_Out_int;
wire	[13:0]FBIO_Out_En_int;

buf	WB_CLK_buf(WB_CLK_int, WB_CLK);
buf	WBs_ACK_buf (WBs_ACK_int, WBs_ACK);
buf	WBs_RD_DAT_buf[31:0] (WBs_RD_DAT_int, WBs_RD_DAT);
buf	SDMA_Req_buf[3:0] (SDMA_Req_int, SDMA_Req);
buf	SDMA_Sreq_buf[3:0] (SDMA_Sreq_int, SDMA_Sreq);
buf	FB_msg_out_buf[3:0] (FB_msg_out_int, FB_msg_out);
buf	FB_Int_Clr_buf[7:0] (FB_Int_Clr_int, FB_Int_Clr);
buf	FB_Busy_buf (FB_Busy_int, FB_Busy);
buf	Sys_PKfb_Clk_buf (Sys_PKfb_Clk_int, Sys_PKfb_Clk);
buf	FB_PKfbData_buf[31:0] (FB_PKfbData_int, FB_PKfbData);
buf	FB_PKfbPush_buf[3:0] (FB_PKfbPush_int, FB_PKfbPush);
buf	Device_ID_buf[15:0] (Device_ID_int, Device_ID);
buf	FBIO_In_En_buf[13:0] (FBIO_In_En_int, FBIO_In_En);
buf	FBIO_Out_buf[13:0] (FBIO_Out_int, FBIO_Out);
buf	FBIO_Out_En_buf[13:0] (FBIO_Out_En_int, FBIO_Out_En);
buf	SPIm_Paddr_buf[15:0] (SPIm_Paddr_int, SPIm_Paddr);
buf	SPIm_PEnable_buf (SPIm_PEnable_int, SPIm_PEnable); 
buf	SPIm_PWdata_buf[31:0] (SPIm_PWdata_int, SPIm_PWdata);
buf	SPIm_PWrite_buf (SPIm_PWrite_int, SPIm_PWrite);
buf	Sys_PSel_buf (Sys_PSel_int, Sys_PSel);
buf FB_PKfbSOF_buf (FB_PKfbSOF_int, FB_PKfbSOF);
buf FB_PKfbEOF_buf (FB_PKfbEOF_int, FB_PKfbEOF);

qlal4s3b_cell_macro inst_qlal4s3b_cell_macro(
						.WB_CLK(WB_CLK_int),
						.WBs_ACK(WBs_ACK_int),
						.WBs_RD_DAT(WBs_RD_DAT_int),
						.WBs_BYTE_STB(WBs_BYTE_STB),
						.WBs_CYC(WBs_CYC),
						.WBs_WE(WBs_WE),
						.WBs_RD(WBs_RD),
						.WBs_STB(WBs_STB),
						.WBs_ADR(WBs_ADR),
						.SDMA_Req(SDMA_Req_int),
						.SDMA_Sreq(SDMA_Sreq_int),
						.SDMA_Done(SDMA_Done),
						.SDMA_Active(SDMA_Active),
						.FB_msg_out(FB_msg_out_int),
						.FB_Int_Clr(FB_Int_Clr_int),		
						.FB_Start(FB_Start),
						.FB_Busy(FB_Busy_int),
						.WB_RST(WB_RST),
						.Sys_PKfb_Rst(Sys_PKfb_Rst),
						.Sys_Clk0(Sys_Clk0),
						.Sys_Clk0_Rst(Sys_Clk0_Rst),
						.Sys_Clk1(Sys_Clk1),
						.Sys_Clk1_Rst(Sys_Clk1_Rst),
						.Sys_Pclk(Sys_Pclk),
						.Sys_Pclk_Rst(Sys_Pclk_Rst),
						.Sys_PKfb_Clk(Sys_PKfb_Clk_int),
						.FB_PKfbData(FB_PKfbData_int),
						.WBs_WR_DAT(WBs_WR_DAT),
						.FB_PKfbPush(FB_PKfbPush_int),
						.FB_PKfbSOF(FB_PKfbSOF_int),
						.FB_PKfbEOF(FB_PKfbEOF_int),
						.Sensor_Int(Sensor_Int),
						.FB_PKfbOverflow(FB_PKfbOverflow),
						.TimeStamp(TimeStamp),
						.Sys_PSel(Sys_PSel_int),
						.SPIm_Paddr(SPIm_Paddr_int),
						.SPIm_PEnable(SPIm_PEnable_int),
						.SPIm_PWrite(SPIm_PWrite_int),
						.SPIm_PWdata(SPIm_PWdata_int),
						.SPIm_PReady(SPIm_PReady),
						.SPIm_PSlvErr(SPIm_PSlvErr),
						.SPIm_Prdata(SPIm_Prdata),
						.Device_ID(Device_ID_int),
						.FBIO_In_En(FBIO_In_En_int),
						.FBIO_Out(FBIO_Out_int),
						.FBIO_Out_En(FBIO_Out_En_int),
						.FBIO_In(FBIO_In),
						.Device_ID_6S(Device_ID_6S), 
						.Device_ID_4S(Device_ID_4S), 
						.SPIm_PWdata_26S(SPIm_PWdata_26S), 
						.SPIm_PWdata_24S(SPIm_PWdata_24S),  
						.SPIm_PWdata_14S(SPIm_PWdata_14S), 
						.SPIm_PWdata_11S(SPIm_PWdata_11S), 
						.SPIm_PWdata_0S(SPIm_PWdata_0S), 
						.SPIm_Paddr_8S(SPIm_Paddr_8S), 
						.SPIm_Paddr_6S(SPIm_Paddr_6S), 
						.FB_PKfbPush_1S(FB_PKfbPush_1S), 
						.FB_PKfbData_31S(FB_PKfbData_31S), 
						.FB_PKfbData_21S(FB_PKfbData_21S),
						.FB_PKfbData_19S(FB_PKfbData_19S),
						.FB_PKfbData_9S(FB_PKfbData_9S),
						.FB_PKfbData_6S(FB_PKfbData_6S),
						.Sys_PKfb_ClkS(Sys_PKfb_ClkS),
						.FB_BusyS(FB_BusyS),
						.WB_CLKS(WB_CLKS),
						.SFBIO(SFBIO)
				);
				
specify
(FB_PKfbPush[3] => FB_PKfbOverflow) = (0,0);
(FB_PKfbPush[2] => FB_PKfbOverflow) = (0,0);
(FB_PKfbPush[1] => FB_PKfbOverflow) = (0,0);
(FB_PKfbPush[0] => FB_PKfbOverflow) = (0,0);
(SPIm_Paddr[11] => SPIm_PReady) = (0,0);
(SPIm_Paddr[10] => SPIm_PReady) = (0,0);
(Sys_PSel => SPIm_PReady) = (0,0);
(SPIm_Paddr[11] => SPIm_PSlvErr) = (0,0);
(SPIm_Paddr[10] => SPIm_PSlvErr) = (0,0);
(Sys_PSel => SPIm_PSlvErr) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[30]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[30]) = (0,0);
(Sys_PSel => SPIm_Prdata[30]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[31]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[31]) = (0,0);
(Sys_PSel => SPIm_Prdata[31]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[22]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[22]) = (0,0);
(Sys_PSel => SPIm_Prdata[22]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[23]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[23]) = (0,0);
(Sys_PSel => SPIm_Prdata[23]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[24]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[24]) = (0,0);
(Sys_PSel => SPIm_Prdata[24]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[25]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[25]) = (0,0);
(Sys_PSel => SPIm_Prdata[25]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[26]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[26]) = (0,0);
(Sys_PSel => SPIm_Prdata[26]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[27]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[27]) = (0,0);
(Sys_PSel => SPIm_Prdata[27]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[28]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[28]) = (0,0);
(Sys_PSel => SPIm_Prdata[28]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[29]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[29]) = (0,0);
(Sys_PSel => SPIm_Prdata[29]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[14]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[14]) = (0,0);
(Sys_PSel => SPIm_Prdata[14]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[15]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[15]) = (0,0);
(Sys_PSel => SPIm_Prdata[15]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[16]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[16]) = (0,0);
(Sys_PSel => SPIm_Prdata[16]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[17]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[17]) = (0,0);
(Sys_PSel => SPIm_Prdata[17]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[18]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[18]) = (0,0);
(Sys_PSel => SPIm_Prdata[18]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[19]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[19]) = (0,0);
(Sys_PSel => SPIm_Prdata[19]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[20]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[20]) = (0,0);
(Sys_PSel => SPIm_Prdata[20]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[21]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[21]) = (0,0);
(Sys_PSel => SPIm_Prdata[21]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[6]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[6]) = (0,0);
(Sys_PSel => SPIm_Prdata[6]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[7]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[7]) = (0,0);
(Sys_PSel => SPIm_Prdata[7]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[8]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[8]) = (0,0);
(Sys_PSel => SPIm_Prdata[8]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[9]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[9]) = (0,0);
(Sys_PSel => SPIm_Prdata[9]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[10]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[10]) = (0,0);
(Sys_PSel => SPIm_Prdata[10]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[11]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[11]) = (0,0);
(Sys_PSel => SPIm_Prdata[11]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[12]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[12]) = (0,0);
(Sys_PSel => SPIm_Prdata[12]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[13]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[13]) = (0,0);
(Sys_PSel => SPIm_Prdata[13]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[0]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[0]) = (0,0);
(Sys_PSel => SPIm_Prdata[0]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[1]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[1]) = (0,0);
(Sys_PSel => SPIm_Prdata[1]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[2]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[2]) = (0,0);
(Sys_PSel => SPIm_Prdata[2]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[3]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[3]) = (0,0);
(Sys_PSel => SPIm_Prdata[3]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[4]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[4]) = (0,0);
(Sys_PSel => SPIm_Prdata[4]) = (0,0);
(SPIm_Paddr[11] => SPIm_Prdata[5]) = (0,0);
(SPIm_Paddr[10] => SPIm_Prdata[5]) = (0,0);
(Sys_PSel => SPIm_Prdata[5]) = (0,0);
(FBIO_In_En[13] => FBIO_In[13]) = (0,0);
(FBIO_In_En[12] => FBIO_In[12]) = (0,0);
(FBIO_In_En[11] => FBIO_In[11]) = (0,0);
(FBIO_In_En[10] => FBIO_In[10]) = (0,0);
(FBIO_In_En[9] => FBIO_In[9]) = (0,0);
(FBIO_In_En[8] => FBIO_In[8]) = (0,0);
(FBIO_In_En[7] => FBIO_In[7]) = (0,0);
(FBIO_In_En[5] => FBIO_In[5]) = (0,0);
(FBIO_In_En[4] => FBIO_In[4]) = (0,0);
(FBIO_In_En[3] => FBIO_In[3]) = (0,0);
(FBIO_In_En[2] => FBIO_In[2]) = (0,0);
(FBIO_In_En[1] => FBIO_In[1]) = (0,0);
(FBIO_In_En[0] => FBIO_In[0]) = (0,0);

endspecify

endmodule

module P_SDIO (IP, IZ, OQI, IE, OE);

input IE, OE, OQI;
output IZ;
inout IP;

assign IZ = IE ? IP : 1'bz;
assign IP = ~OE ? OQI : 1'bz;

specify

if ( IE == 1'b1 ) (IP => IZ) = (0,0);
if ( OE == 1'b0 ) (OQI => IP) = (0,0);

(IE => IP) = (0,0,0,0,0,0);
(OE => IP) = (0,0,0,0,0,0);

endspecify

endmodule
