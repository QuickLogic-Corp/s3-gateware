

module decimation_filter_3to1 (
);


