
`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE0_PR0_WSA0_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A2_b0, posedge CLK2, "");
      $hold(posedge CLK2, A2_b0, "");
      $setup(A2_b1, posedge CLK2, "");
      $hold(posedge CLK2, A2_b1, "");
      $setup(A2_b2, posedge CLK2, "");
      $hold(posedge CLK2, A2_b2, "");
      $setup(A2_b3, posedge CLK2, "");
      $hold(posedge CLK2, A2_b3, "");
      $setup(A2_b4, posedge CLK2, "");
      $hold(posedge CLK2, A2_b4, "");
      $setup(A2_b5, posedge CLK2, "");
      $hold(posedge CLK2, A2_b5, "");
      $setup(A2_b6, posedge CLK2, "");
      $hold(posedge CLK2, A2_b6, "");
      $setup(A2_b7, posedge CLK2, "");
      $hold(posedge CLK2, A2_b7, "");
      $setup(A2_b8, posedge CLK2, "");
      $hold(posedge CLK2, A2_b8, "");
      $setup(A2_b9, posedge CLK2, "");
      $hold(posedge CLK2, A2_b9, "");
      $setup(A2_b10, posedge CLK2, "");
      $hold(posedge CLK2, A2_b10, "");
      $setup(WEN1_b0, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b0, "");
      $setup(WEN1_b1, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b1, "");
      $setup(A1_b0, posedge CLK1, "");
      $hold(posedge CLK1, A1_b0, "");
      $setup(A1_b1, posedge CLK1, "");
      $hold(posedge CLK1, A1_b1, "");
      $setup(A1_b2, posedge CLK1, "");
      $hold(posedge CLK1, A1_b2, "");
      $setup(A1_b3, posedge CLK1, "");
      $hold(posedge CLK1, A1_b3, "");
      $setup(A1_b4, posedge CLK1, "");
      $hold(posedge CLK1, A1_b4, "");
      $setup(A1_b5, posedge CLK1, "");
      $hold(posedge CLK1, A1_b5, "");
      $setup(A1_b6, posedge CLK1, "");
      $hold(posedge CLK1, A1_b6, "");
      $setup(A1_b7, posedge CLK1, "");
      $hold(posedge CLK1, A1_b7, "");
      $setup(A1_b8, posedge CLK1, "");
      $hold(posedge CLK1, A1_b8, "");
      $setup(A1_b9, posedge CLK1, "");
      $hold(posedge CLK1, A1_b9, "");
      $setup(A1_b10, posedge CLK1, "");
      $hold(posedge CLK1, A1_b10, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE0_PR0_WSA0_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A2_b0, posedge CLK2, "");
      $hold(posedge CLK2, A2_b0, "");
      $setup(A2_b1, posedge CLK2, "");
      $hold(posedge CLK2, A2_b1, "");
      $setup(A2_b2, posedge CLK2, "");
      $hold(posedge CLK2, A2_b2, "");
      $setup(A2_b3, posedge CLK2, "");
      $hold(posedge CLK2, A2_b3, "");
      $setup(A2_b4, posedge CLK2, "");
      $hold(posedge CLK2, A2_b4, "");
      $setup(A2_b5, posedge CLK2, "");
      $hold(posedge CLK2, A2_b5, "");
      $setup(A2_b6, posedge CLK2, "");
      $hold(posedge CLK2, A2_b6, "");
      $setup(A2_b7, posedge CLK2, "");
      $hold(posedge CLK2, A2_b7, "");
      $setup(A2_b8, posedge CLK2, "");
      $hold(posedge CLK2, A2_b8, "");
      $setup(A2_b9, posedge CLK2, "");
      $hold(posedge CLK2, A2_b9, "");
      $setup(A2_b10, posedge CLK2, "");
      $hold(posedge CLK2, A2_b10, "");
      $setup(WEN1_b0, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b0, "");
      $setup(WEN1_b1, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b1, "");
      $setup(A1_b0, posedge CLK1, "");
      $hold(posedge CLK1, A1_b0, "");
      $setup(A1_b1, posedge CLK1, "");
      $hold(posedge CLK1, A1_b1, "");
      $setup(A1_b2, posedge CLK1, "");
      $hold(posedge CLK1, A1_b2, "");
      $setup(A1_b3, posedge CLK1, "");
      $hold(posedge CLK1, A1_b3, "");
      $setup(A1_b4, posedge CLK1, "");
      $hold(posedge CLK1, A1_b4, "");
      $setup(A1_b5, posedge CLK1, "");
      $hold(posedge CLK1, A1_b5, "");
      $setup(A1_b6, posedge CLK1, "");
      $hold(posedge CLK1, A1_b6, "");
      $setup(A1_b7, posedge CLK1, "");
      $hold(posedge CLK1, A1_b7, "");
      $setup(A1_b8, posedge CLK1, "");
      $hold(posedge CLK1, A1_b8, "");
      $setup(A1_b9, posedge CLK1, "");
      $hold(posedge CLK1, A1_b9, "");
      $setup(A1_b10, posedge CLK1, "");
      $hold(posedge CLK1, A1_b10, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE0_PR0_WSA1_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A2_b0, posedge CLK2, "");
      $hold(posedge CLK2, A2_b0, "");
      $setup(A2_b1, posedge CLK2, "");
      $hold(posedge CLK2, A2_b1, "");
      $setup(A2_b2, posedge CLK2, "");
      $hold(posedge CLK2, A2_b2, "");
      $setup(A2_b3, posedge CLK2, "");
      $hold(posedge CLK2, A2_b3, "");
      $setup(A2_b4, posedge CLK2, "");
      $hold(posedge CLK2, A2_b4, "");
      $setup(A2_b5, posedge CLK2, "");
      $hold(posedge CLK2, A2_b5, "");
      $setup(A2_b6, posedge CLK2, "");
      $hold(posedge CLK2, A2_b6, "");
      $setup(A2_b7, posedge CLK2, "");
      $hold(posedge CLK2, A2_b7, "");
      $setup(A2_b8, posedge CLK2, "");
      $hold(posedge CLK2, A2_b8, "");
      $setup(A2_b9, posedge CLK2, "");
      $hold(posedge CLK2, A2_b9, "");
      $setup(A2_b10, posedge CLK2, "");
      $hold(posedge CLK2, A2_b10, "");
      $setup(WEN1_b0, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b0, "");
      $setup(WEN1_b1, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b1, "");
      $setup(A1_b0, posedge CLK1, "");
      $hold(posedge CLK1, A1_b0, "");
      $setup(A1_b1, posedge CLK1, "");
      $hold(posedge CLK1, A1_b1, "");
      $setup(A1_b2, posedge CLK1, "");
      $hold(posedge CLK1, A1_b2, "");
      $setup(A1_b3, posedge CLK1, "");
      $hold(posedge CLK1, A1_b3, "");
      $setup(A1_b4, posedge CLK1, "");
      $hold(posedge CLK1, A1_b4, "");
      $setup(A1_b5, posedge CLK1, "");
      $hold(posedge CLK1, A1_b5, "");
      $setup(A1_b6, posedge CLK1, "");
      $hold(posedge CLK1, A1_b6, "");
      $setup(A1_b7, posedge CLK1, "");
      $hold(posedge CLK1, A1_b7, "");
      $setup(A1_b8, posedge CLK1, "");
      $hold(posedge CLK1, A1_b8, "");
      $setup(A1_b9, posedge CLK1, "");
      $hold(posedge CLK1, A1_b9, "");
      $setup(A1_b10, posedge CLK1, "");
      $hold(posedge CLK1, A1_b10, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE0_PR0_WSA1_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A2_b0, posedge CLK2, "");
      $hold(posedge CLK2, A2_b0, "");
      $setup(A2_b1, posedge CLK2, "");
      $hold(posedge CLK2, A2_b1, "");
      $setup(A2_b2, posedge CLK2, "");
      $hold(posedge CLK2, A2_b2, "");
      $setup(A2_b3, posedge CLK2, "");
      $hold(posedge CLK2, A2_b3, "");
      $setup(A2_b4, posedge CLK2, "");
      $hold(posedge CLK2, A2_b4, "");
      $setup(A2_b5, posedge CLK2, "");
      $hold(posedge CLK2, A2_b5, "");
      $setup(A2_b6, posedge CLK2, "");
      $hold(posedge CLK2, A2_b6, "");
      $setup(A2_b7, posedge CLK2, "");
      $hold(posedge CLK2, A2_b7, "");
      $setup(A2_b8, posedge CLK2, "");
      $hold(posedge CLK2, A2_b8, "");
      $setup(A2_b9, posedge CLK2, "");
      $hold(posedge CLK2, A2_b9, "");
      $setup(A2_b10, posedge CLK2, "");
      $hold(posedge CLK2, A2_b10, "");
      $setup(WEN1_b0, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b0, "");
      $setup(WEN1_b1, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b1, "");
      $setup(A1_b0, posedge CLK1, "");
      $hold(posedge CLK1, A1_b0, "");
      $setup(A1_b1, posedge CLK1, "");
      $hold(posedge CLK1, A1_b1, "");
      $setup(A1_b2, posedge CLK1, "");
      $hold(posedge CLK1, A1_b2, "");
      $setup(A1_b3, posedge CLK1, "");
      $hold(posedge CLK1, A1_b3, "");
      $setup(A1_b4, posedge CLK1, "");
      $hold(posedge CLK1, A1_b4, "");
      $setup(A1_b5, posedge CLK1, "");
      $hold(posedge CLK1, A1_b5, "");
      $setup(A1_b6, posedge CLK1, "");
      $hold(posedge CLK1, A1_b6, "");
      $setup(A1_b7, posedge CLK1, "");
      $hold(posedge CLK1, A1_b7, "");
      $setup(A1_b8, posedge CLK1, "");
      $hold(posedge CLK1, A1_b8, "");
      $setup(A1_b9, posedge CLK1, "");
      $hold(posedge CLK1, A1_b9, "");
      $setup(A1_b10, posedge CLK1, "");
      $hold(posedge CLK1, A1_b10, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE0_PR1_WSA0_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A2_b0, posedge CLK2, "");
      $hold(posedge CLK2, A2_b0, "");
      $setup(A2_b1, posedge CLK2, "");
      $hold(posedge CLK2, A2_b1, "");
      $setup(A2_b2, posedge CLK2, "");
      $hold(posedge CLK2, A2_b2, "");
      $setup(A2_b3, posedge CLK2, "");
      $hold(posedge CLK2, A2_b3, "");
      $setup(A2_b4, posedge CLK2, "");
      $hold(posedge CLK2, A2_b4, "");
      $setup(A2_b5, posedge CLK2, "");
      $hold(posedge CLK2, A2_b5, "");
      $setup(A2_b6, posedge CLK2, "");
      $hold(posedge CLK2, A2_b6, "");
      $setup(A2_b7, posedge CLK2, "");
      $hold(posedge CLK2, A2_b7, "");
      $setup(A2_b8, posedge CLK2, "");
      $hold(posedge CLK2, A2_b8, "");
      $setup(A2_b9, posedge CLK2, "");
      $hold(posedge CLK2, A2_b9, "");
      $setup(A2_b10, posedge CLK2, "");
      $hold(posedge CLK2, A2_b10, "");
      $setup(WEN1_b0, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b0, "");
      $setup(WEN1_b1, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b1, "");
      $setup(A1_b0, posedge CLK1, "");
      $hold(posedge CLK1, A1_b0, "");
      $setup(A1_b1, posedge CLK1, "");
      $hold(posedge CLK1, A1_b1, "");
      $setup(A1_b2, posedge CLK1, "");
      $hold(posedge CLK1, A1_b2, "");
      $setup(A1_b3, posedge CLK1, "");
      $hold(posedge CLK1, A1_b3, "");
      $setup(A1_b4, posedge CLK1, "");
      $hold(posedge CLK1, A1_b4, "");
      $setup(A1_b5, posedge CLK1, "");
      $hold(posedge CLK1, A1_b5, "");
      $setup(A1_b6, posedge CLK1, "");
      $hold(posedge CLK1, A1_b6, "");
      $setup(A1_b7, posedge CLK1, "");
      $hold(posedge CLK1, A1_b7, "");
      $setup(A1_b8, posedge CLK1, "");
      $hold(posedge CLK1, A1_b8, "");
      $setup(A1_b9, posedge CLK1, "");
      $hold(posedge CLK1, A1_b9, "");
      $setup(A1_b10, posedge CLK1, "");
      $hold(posedge CLK1, A1_b10, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE0_PR1_WSA0_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A2_b0, posedge CLK2, "");
      $hold(posedge CLK2, A2_b0, "");
      $setup(A2_b1, posedge CLK2, "");
      $hold(posedge CLK2, A2_b1, "");
      $setup(A2_b2, posedge CLK2, "");
      $hold(posedge CLK2, A2_b2, "");
      $setup(A2_b3, posedge CLK2, "");
      $hold(posedge CLK2, A2_b3, "");
      $setup(A2_b4, posedge CLK2, "");
      $hold(posedge CLK2, A2_b4, "");
      $setup(A2_b5, posedge CLK2, "");
      $hold(posedge CLK2, A2_b5, "");
      $setup(A2_b6, posedge CLK2, "");
      $hold(posedge CLK2, A2_b6, "");
      $setup(A2_b7, posedge CLK2, "");
      $hold(posedge CLK2, A2_b7, "");
      $setup(A2_b8, posedge CLK2, "");
      $hold(posedge CLK2, A2_b8, "");
      $setup(A2_b9, posedge CLK2, "");
      $hold(posedge CLK2, A2_b9, "");
      $setup(A2_b10, posedge CLK2, "");
      $hold(posedge CLK2, A2_b10, "");
      $setup(WEN1_b0, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b0, "");
      $setup(WEN1_b1, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b1, "");
      $setup(A1_b0, posedge CLK1, "");
      $hold(posedge CLK1, A1_b0, "");
      $setup(A1_b1, posedge CLK1, "");
      $hold(posedge CLK1, A1_b1, "");
      $setup(A1_b2, posedge CLK1, "");
      $hold(posedge CLK1, A1_b2, "");
      $setup(A1_b3, posedge CLK1, "");
      $hold(posedge CLK1, A1_b3, "");
      $setup(A1_b4, posedge CLK1, "");
      $hold(posedge CLK1, A1_b4, "");
      $setup(A1_b5, posedge CLK1, "");
      $hold(posedge CLK1, A1_b5, "");
      $setup(A1_b6, posedge CLK1, "");
      $hold(posedge CLK1, A1_b6, "");
      $setup(A1_b7, posedge CLK1, "");
      $hold(posedge CLK1, A1_b7, "");
      $setup(A1_b8, posedge CLK1, "");
      $hold(posedge CLK1, A1_b8, "");
      $setup(A1_b9, posedge CLK1, "");
      $hold(posedge CLK1, A1_b9, "");
      $setup(A1_b10, posedge CLK1, "");
      $hold(posedge CLK1, A1_b10, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE0_PR1_WSA1_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A2_b0, posedge CLK2, "");
      $hold(posedge CLK2, A2_b0, "");
      $setup(A2_b1, posedge CLK2, "");
      $hold(posedge CLK2, A2_b1, "");
      $setup(A2_b2, posedge CLK2, "");
      $hold(posedge CLK2, A2_b2, "");
      $setup(A2_b3, posedge CLK2, "");
      $hold(posedge CLK2, A2_b3, "");
      $setup(A2_b4, posedge CLK2, "");
      $hold(posedge CLK2, A2_b4, "");
      $setup(A2_b5, posedge CLK2, "");
      $hold(posedge CLK2, A2_b5, "");
      $setup(A2_b6, posedge CLK2, "");
      $hold(posedge CLK2, A2_b6, "");
      $setup(A2_b7, posedge CLK2, "");
      $hold(posedge CLK2, A2_b7, "");
      $setup(A2_b8, posedge CLK2, "");
      $hold(posedge CLK2, A2_b8, "");
      $setup(A2_b9, posedge CLK2, "");
      $hold(posedge CLK2, A2_b9, "");
      $setup(A2_b10, posedge CLK2, "");
      $hold(posedge CLK2, A2_b10, "");
      $setup(WEN1_b0, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b0, "");
      $setup(WEN1_b1, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b1, "");
      $setup(A1_b0, posedge CLK1, "");
      $hold(posedge CLK1, A1_b0, "");
      $setup(A1_b1, posedge CLK1, "");
      $hold(posedge CLK1, A1_b1, "");
      $setup(A1_b2, posedge CLK1, "");
      $hold(posedge CLK1, A1_b2, "");
      $setup(A1_b3, posedge CLK1, "");
      $hold(posedge CLK1, A1_b3, "");
      $setup(A1_b4, posedge CLK1, "");
      $hold(posedge CLK1, A1_b4, "");
      $setup(A1_b5, posedge CLK1, "");
      $hold(posedge CLK1, A1_b5, "");
      $setup(A1_b6, posedge CLK1, "");
      $hold(posedge CLK1, A1_b6, "");
      $setup(A1_b7, posedge CLK1, "");
      $hold(posedge CLK1, A1_b7, "");
      $setup(A1_b8, posedge CLK1, "");
      $hold(posedge CLK1, A1_b8, "");
      $setup(A1_b9, posedge CLK1, "");
      $hold(posedge CLK1, A1_b9, "");
      $setup(A1_b10, posedge CLK1, "");
      $hold(posedge CLK1, A1_b10, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE0_PR1_WSA1_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A2_b0, posedge CLK2, "");
      $hold(posedge CLK2, A2_b0, "");
      $setup(A2_b1, posedge CLK2, "");
      $hold(posedge CLK2, A2_b1, "");
      $setup(A2_b2, posedge CLK2, "");
      $hold(posedge CLK2, A2_b2, "");
      $setup(A2_b3, posedge CLK2, "");
      $hold(posedge CLK2, A2_b3, "");
      $setup(A2_b4, posedge CLK2, "");
      $hold(posedge CLK2, A2_b4, "");
      $setup(A2_b5, posedge CLK2, "");
      $hold(posedge CLK2, A2_b5, "");
      $setup(A2_b6, posedge CLK2, "");
      $hold(posedge CLK2, A2_b6, "");
      $setup(A2_b7, posedge CLK2, "");
      $hold(posedge CLK2, A2_b7, "");
      $setup(A2_b8, posedge CLK2, "");
      $hold(posedge CLK2, A2_b8, "");
      $setup(A2_b9, posedge CLK2, "");
      $hold(posedge CLK2, A2_b9, "");
      $setup(A2_b10, posedge CLK2, "");
      $hold(posedge CLK2, A2_b10, "");
      $setup(WEN1_b0, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b0, "");
      $setup(WEN1_b1, posedge CLK1, "");
      $hold(posedge CLK1, WEN1_b1, "");
      $setup(A1_b0, posedge CLK1, "");
      $hold(posedge CLK1, A1_b0, "");
      $setup(A1_b1, posedge CLK1, "");
      $hold(posedge CLK1, A1_b1, "");
      $setup(A1_b2, posedge CLK1, "");
      $hold(posedge CLK1, A1_b2, "");
      $setup(A1_b3, posedge CLK1, "");
      $hold(posedge CLK1, A1_b3, "");
      $setup(A1_b4, posedge CLK1, "");
      $hold(posedge CLK1, A1_b4, "");
      $setup(A1_b5, posedge CLK1, "");
      $hold(posedge CLK1, A1_b5, "");
      $setup(A1_b6, posedge CLK1, "");
      $hold(posedge CLK1, A1_b6, "");
      $setup(A1_b7, posedge CLK1, "");
      $hold(posedge CLK1, A1_b7, "");
      $setup(A1_b8, posedge CLK1, "");
      $hold(posedge CLK1, A1_b8, "");
      $setup(A1_b9, posedge CLK1, "");
      $hold(posedge CLK1, A1_b9, "");
      $setup(A1_b10, posedge CLK1, "");
      $hold(posedge CLK1, A1_b10, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D0_PR0_WSA0_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>Almost_Full)="";
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
      (CLK2*>Almost_Empty)="";
      (CLK1*>PUSH_FLAG_b0)="";
      (CLK1*>PUSH_FLAG_b1)="";
      (CLK1*>PUSH_FLAG_b2)="";
      (CLK1*>PUSH_FLAG_b3)="";
      (CLK2*>POP_FLAG_b0)="";
      (CLK2*>POP_FLAG_b1)="";
      (CLK2*>POP_FLAG_b2)="";
      (CLK2*>POP_FLAG_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D0_PR0_WSA0_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>Almost_Full)="";
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
      (CLK2*>Almost_Empty)="";
      (CLK1*>PUSH_FLAG_b0)="";
      (CLK1*>PUSH_FLAG_b1)="";
      (CLK1*>PUSH_FLAG_b2)="";
      (CLK1*>PUSH_FLAG_b3)="";
      (CLK2*>POP_FLAG_b0)="";
      (CLK2*>POP_FLAG_b1)="";
      (CLK2*>POP_FLAG_b2)="";
      (CLK2*>POP_FLAG_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D0_PR0_WSA1_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>Almost_Full)="";
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
      (CLK2*>Almost_Empty)="";
      (CLK1*>PUSH_FLAG_b0)="";
      (CLK1*>PUSH_FLAG_b1)="";
      (CLK1*>PUSH_FLAG_b2)="";
      (CLK1*>PUSH_FLAG_b3)="";
      (CLK2*>POP_FLAG_b0)="";
      (CLK2*>POP_FLAG_b1)="";
      (CLK2*>POP_FLAG_b2)="";
      (CLK2*>POP_FLAG_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D0_PR0_WSA1_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>Almost_Full)="";
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
      (CLK2*>Almost_Empty)="";
      (CLK1*>PUSH_FLAG_b0)="";
      (CLK1*>PUSH_FLAG_b1)="";
      (CLK1*>PUSH_FLAG_b2)="";
      (CLK1*>PUSH_FLAG_b3)="";
      (CLK2*>POP_FLAG_b0)="";
      (CLK2*>POP_FLAG_b1)="";
      (CLK2*>POP_FLAG_b2)="";
      (CLK2*>POP_FLAG_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D0_PR1_WSA0_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>Almost_Full)="";
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
      (CLK2*>Almost_Empty)="";
      (CLK1*>PUSH_FLAG_b0)="";
      (CLK1*>PUSH_FLAG_b1)="";
      (CLK1*>PUSH_FLAG_b2)="";
      (CLK1*>PUSH_FLAG_b3)="";
      (CLK2*>POP_FLAG_b0)="";
      (CLK2*>POP_FLAG_b1)="";
      (CLK2*>POP_FLAG_b2)="";
      (CLK2*>POP_FLAG_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D0_PR1_WSA0_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>Almost_Full)="";
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
      (CLK2*>Almost_Empty)="";
      (CLK1*>PUSH_FLAG_b0)="";
      (CLK1*>PUSH_FLAG_b1)="";
      (CLK1*>PUSH_FLAG_b2)="";
      (CLK1*>PUSH_FLAG_b3)="";
      (CLK2*>POP_FLAG_b0)="";
      (CLK2*>POP_FLAG_b1)="";
      (CLK2*>POP_FLAG_b2)="";
      (CLK2*>POP_FLAG_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D0_PR1_WSA1_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>Almost_Full)="";
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
      (CLK2*>Almost_Empty)="";
      (CLK1*>PUSH_FLAG_b0)="";
      (CLK1*>PUSH_FLAG_b1)="";
      (CLK1*>PUSH_FLAG_b2)="";
      (CLK1*>PUSH_FLAG_b3)="";
      (CLK2*>POP_FLAG_b0)="";
      (CLK2*>POP_FLAG_b1)="";
      (CLK2*>POP_FLAG_b2)="";
      (CLK2*>POP_FLAG_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D0_PR1_WSA1_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         TEST1B,
  input         PIPELINE_RD,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         WEN1_b0,
  input         WEN1_b1,
  input         LS,
  input         SD_RB1,
  input         CS1,
  input         TEST1A,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        Almost_Full,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Empty,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK1, "");
      $hold(posedge CLK1, WD_b0, "");
      $setup(WD_b1, posedge CLK1, "");
      $hold(posedge CLK1, WD_b1, "");
      $setup(WD_b2, posedge CLK1, "");
      $hold(posedge CLK1, WD_b2, "");
      $setup(WD_b3, posedge CLK1, "");
      $hold(posedge CLK1, WD_b3, "");
      $setup(WD_b4, posedge CLK1, "");
      $hold(posedge CLK1, WD_b4, "");
      $setup(WD_b5, posedge CLK1, "");
      $hold(posedge CLK1, WD_b5, "");
      $setup(WD_b6, posedge CLK1, "");
      $hold(posedge CLK1, WD_b6, "");
      $setup(WD_b7, posedge CLK1, "");
      $hold(posedge CLK1, WD_b7, "");
      $setup(WD_b8, posedge CLK1, "");
      $hold(posedge CLK1, WD_b8, "");
      $setup(WD_b9, posedge CLK1, "");
      $hold(posedge CLK1, WD_b9, "");
      $setup(WD_b10, posedge CLK1, "");
      $hold(posedge CLK1, WD_b10, "");
      $setup(WD_b11, posedge CLK1, "");
      $hold(posedge CLK1, WD_b11, "");
      $setup(WD_b12, posedge CLK1, "");
      $hold(posedge CLK1, WD_b12, "");
      $setup(WD_b13, posedge CLK1, "");
      $hold(posedge CLK1, WD_b13, "");
      $setup(WD_b14, posedge CLK1, "");
      $hold(posedge CLK1, WD_b14, "");
      $setup(WD_b15, posedge CLK1, "");
      $hold(posedge CLK1, WD_b15, "");
      $setup(WD_b16, posedge CLK1, "");
      $hold(posedge CLK1, WD_b16, "");
      $setup(WD_b17, posedge CLK1, "");
      $hold(posedge CLK1, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>Almost_Full)="";
      (CLK2*>RD_b0)="";
      (CLK2*>RD_b1)="";
      (CLK2*>RD_b2)="";
      (CLK2*>RD_b3)="";
      (CLK2*>RD_b4)="";
      (CLK2*>RD_b5)="";
      (CLK2*>RD_b6)="";
      (CLK2*>RD_b7)="";
      (CLK2*>RD_b8)="";
      (CLK2*>RD_b9)="";
      (CLK2*>RD_b10)="";
      (CLK2*>RD_b11)="";
      (CLK2*>RD_b12)="";
      (CLK2*>RD_b13)="";
      (CLK2*>RD_b14)="";
      (CLK2*>RD_b15)="";
      (CLK2*>RD_b16)="";
      (CLK2*>RD_b17)="";
      (CLK2*>Almost_Empty)="";
      (CLK1*>PUSH_FLAG_b0)="";
      (CLK1*>PUSH_FLAG_b1)="";
      (CLK1*>PUSH_FLAG_b2)="";
      (CLK1*>PUSH_FLAG_b3)="";
      (CLK2*>POP_FLAG_b0)="";
      (CLK2*>POP_FLAG_b1)="";
      (CLK2*>POP_FLAG_b2)="";
      (CLK2*>POP_FLAG_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .P1_0(P1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .Almost_Full_0(Almost_Full),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Empty_0(Almost_Empty),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D1_PR0_WSA0_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         TEST1B,
  input         PIPELINE_RD,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         LS,
  input         SD_RB1,
  input         TEST1A,
  input         CS1,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_b0,
  input         WEN1_b1,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Full,
  output        Almost_Empty
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK2, "");
      $hold(posedge CLK2, WD_b0, "");
      $setup(WD_b1, posedge CLK2, "");
      $hold(posedge CLK2, WD_b1, "");
      $setup(WD_b2, posedge CLK2, "");
      $hold(posedge CLK2, WD_b2, "");
      $setup(WD_b3, posedge CLK2, "");
      $hold(posedge CLK2, WD_b3, "");
      $setup(WD_b4, posedge CLK2, "");
      $hold(posedge CLK2, WD_b4, "");
      $setup(WD_b5, posedge CLK2, "");
      $hold(posedge CLK2, WD_b5, "");
      $setup(WD_b6, posedge CLK2, "");
      $hold(posedge CLK2, WD_b6, "");
      $setup(WD_b7, posedge CLK2, "");
      $hold(posedge CLK2, WD_b7, "");
      $setup(WD_b8, posedge CLK2, "");
      $hold(posedge CLK2, WD_b8, "");
      $setup(WD_b9, posedge CLK2, "");
      $hold(posedge CLK2, WD_b9, "");
      $setup(WD_b10, posedge CLK2, "");
      $hold(posedge CLK2, WD_b10, "");
      $setup(WD_b11, posedge CLK2, "");
      $hold(posedge CLK2, WD_b11, "");
      $setup(WD_b12, posedge CLK2, "");
      $hold(posedge CLK2, WD_b12, "");
      $setup(WD_b13, posedge CLK2, "");
      $hold(posedge CLK2, WD_b13, "");
      $setup(WD_b14, posedge CLK2, "");
      $hold(posedge CLK2, WD_b14, "");
      $setup(WD_b15, posedge CLK2, "");
      $hold(posedge CLK2, WD_b15, "");
      $setup(WD_b16, posedge CLK2, "");
      $hold(posedge CLK2, WD_b16, "");
      $setup(WD_b17, posedge CLK2, "");
      $hold(posedge CLK2, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>POP_FLAG_b0)="";
      (CLK1*>POP_FLAG_b1)="";
      (CLK1*>POP_FLAG_b2)="";
      (CLK1*>POP_FLAG_b3)="";
      (CLK2*>PUSH_FLAG_b0)="";
      (CLK2*>PUSH_FLAG_b1)="";
      (CLK2*>PUSH_FLAG_b2)="";
      (CLK2*>PUSH_FLAG_b3)="";
      (CLK1*>RD_b0)="";
      (CLK1*>RD_b1)="";
      (CLK1*>RD_b2)="";
      (CLK1*>RD_b3)="";
      (CLK1*>RD_b4)="";
      (CLK1*>RD_b5)="";
      (CLK1*>RD_b6)="";
      (CLK1*>RD_b7)="";
      (CLK1*>RD_b8)="";
      (CLK1*>RD_b9)="";
      (CLK1*>RD_b10)="";
      (CLK1*>RD_b11)="";
      (CLK1*>RD_b12)="";
      (CLK1*>RD_b13)="";
      (CLK1*>RD_b14)="";
      (CLK1*>RD_b15)="";
      (CLK1*>RD_b16)="";
      (CLK1*>RD_b17)="";
      (CLK2*>Almost_Full)="";
      (CLK1*>Almost_Empty)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .P1_0(P1),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Full_0(Almost_Full),
      .Almost_Empty_0(Almost_Empty));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D1_PR0_WSA0_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         TEST1B,
  input         PIPELINE_RD,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         LS,
  input         SD_RB1,
  input         TEST1A,
  input         CS1,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_b0,
  input         WEN1_b1,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Full,
  output        Almost_Empty
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK2, "");
      $hold(posedge CLK2, WD_b0, "");
      $setup(WD_b1, posedge CLK2, "");
      $hold(posedge CLK2, WD_b1, "");
      $setup(WD_b2, posedge CLK2, "");
      $hold(posedge CLK2, WD_b2, "");
      $setup(WD_b3, posedge CLK2, "");
      $hold(posedge CLK2, WD_b3, "");
      $setup(WD_b4, posedge CLK2, "");
      $hold(posedge CLK2, WD_b4, "");
      $setup(WD_b5, posedge CLK2, "");
      $hold(posedge CLK2, WD_b5, "");
      $setup(WD_b6, posedge CLK2, "");
      $hold(posedge CLK2, WD_b6, "");
      $setup(WD_b7, posedge CLK2, "");
      $hold(posedge CLK2, WD_b7, "");
      $setup(WD_b8, posedge CLK2, "");
      $hold(posedge CLK2, WD_b8, "");
      $setup(WD_b9, posedge CLK2, "");
      $hold(posedge CLK2, WD_b9, "");
      $setup(WD_b10, posedge CLK2, "");
      $hold(posedge CLK2, WD_b10, "");
      $setup(WD_b11, posedge CLK2, "");
      $hold(posedge CLK2, WD_b11, "");
      $setup(WD_b12, posedge CLK2, "");
      $hold(posedge CLK2, WD_b12, "");
      $setup(WD_b13, posedge CLK2, "");
      $hold(posedge CLK2, WD_b13, "");
      $setup(WD_b14, posedge CLK2, "");
      $hold(posedge CLK2, WD_b14, "");
      $setup(WD_b15, posedge CLK2, "");
      $hold(posedge CLK2, WD_b15, "");
      $setup(WD_b16, posedge CLK2, "");
      $hold(posedge CLK2, WD_b16, "");
      $setup(WD_b17, posedge CLK2, "");
      $hold(posedge CLK2, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>POP_FLAG_b0)="";
      (CLK1*>POP_FLAG_b1)="";
      (CLK1*>POP_FLAG_b2)="";
      (CLK1*>POP_FLAG_b3)="";
      (CLK2*>PUSH_FLAG_b0)="";
      (CLK2*>PUSH_FLAG_b1)="";
      (CLK2*>PUSH_FLAG_b2)="";
      (CLK2*>PUSH_FLAG_b3)="";
      (CLK1*>RD_b0)="";
      (CLK1*>RD_b1)="";
      (CLK1*>RD_b2)="";
      (CLK1*>RD_b3)="";
      (CLK1*>RD_b4)="";
      (CLK1*>RD_b5)="";
      (CLK1*>RD_b6)="";
      (CLK1*>RD_b7)="";
      (CLK1*>RD_b8)="";
      (CLK1*>RD_b9)="";
      (CLK1*>RD_b10)="";
      (CLK1*>RD_b11)="";
      (CLK1*>RD_b12)="";
      (CLK1*>RD_b13)="";
      (CLK1*>RD_b14)="";
      (CLK1*>RD_b15)="";
      (CLK1*>RD_b16)="";
      (CLK1*>RD_b17)="";
      (CLK2*>Almost_Full)="";
      (CLK1*>Almost_Empty)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .P1_0(P1),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Full_0(Almost_Full),
      .Almost_Empty_0(Almost_Empty));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D1_PR0_WSA1_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         TEST1B,
  input         PIPELINE_RD,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         LS,
  input         SD_RB1,
  input         TEST1A,
  input         CS1,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_b0,
  input         WEN1_b1,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Full,
  output        Almost_Empty
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK2, "");
      $hold(posedge CLK2, WD_b0, "");
      $setup(WD_b1, posedge CLK2, "");
      $hold(posedge CLK2, WD_b1, "");
      $setup(WD_b2, posedge CLK2, "");
      $hold(posedge CLK2, WD_b2, "");
      $setup(WD_b3, posedge CLK2, "");
      $hold(posedge CLK2, WD_b3, "");
      $setup(WD_b4, posedge CLK2, "");
      $hold(posedge CLK2, WD_b4, "");
      $setup(WD_b5, posedge CLK2, "");
      $hold(posedge CLK2, WD_b5, "");
      $setup(WD_b6, posedge CLK2, "");
      $hold(posedge CLK2, WD_b6, "");
      $setup(WD_b7, posedge CLK2, "");
      $hold(posedge CLK2, WD_b7, "");
      $setup(WD_b8, posedge CLK2, "");
      $hold(posedge CLK2, WD_b8, "");
      $setup(WD_b9, posedge CLK2, "");
      $hold(posedge CLK2, WD_b9, "");
      $setup(WD_b10, posedge CLK2, "");
      $hold(posedge CLK2, WD_b10, "");
      $setup(WD_b11, posedge CLK2, "");
      $hold(posedge CLK2, WD_b11, "");
      $setup(WD_b12, posedge CLK2, "");
      $hold(posedge CLK2, WD_b12, "");
      $setup(WD_b13, posedge CLK2, "");
      $hold(posedge CLK2, WD_b13, "");
      $setup(WD_b14, posedge CLK2, "");
      $hold(posedge CLK2, WD_b14, "");
      $setup(WD_b15, posedge CLK2, "");
      $hold(posedge CLK2, WD_b15, "");
      $setup(WD_b16, posedge CLK2, "");
      $hold(posedge CLK2, WD_b16, "");
      $setup(WD_b17, posedge CLK2, "");
      $hold(posedge CLK2, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>POP_FLAG_b0)="";
      (CLK1*>POP_FLAG_b1)="";
      (CLK1*>POP_FLAG_b2)="";
      (CLK1*>POP_FLAG_b3)="";
      (CLK2*>PUSH_FLAG_b0)="";
      (CLK2*>PUSH_FLAG_b1)="";
      (CLK2*>PUSH_FLAG_b2)="";
      (CLK2*>PUSH_FLAG_b3)="";
      (CLK1*>RD_b0)="";
      (CLK1*>RD_b1)="";
      (CLK1*>RD_b2)="";
      (CLK1*>RD_b3)="";
      (CLK1*>RD_b4)="";
      (CLK1*>RD_b5)="";
      (CLK1*>RD_b6)="";
      (CLK1*>RD_b7)="";
      (CLK1*>RD_b8)="";
      (CLK1*>RD_b9)="";
      (CLK1*>RD_b10)="";
      (CLK1*>RD_b11)="";
      (CLK1*>RD_b12)="";
      (CLK1*>RD_b13)="";
      (CLK1*>RD_b14)="";
      (CLK1*>RD_b15)="";
      (CLK1*>RD_b16)="";
      (CLK1*>RD_b17)="";
      (CLK2*>Almost_Full)="";
      (CLK1*>Almost_Empty)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .P1_0(P1),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Full_0(Almost_Full),
      .Almost_Empty_0(Almost_Empty));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D1_PR0_WSA1_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         TEST1B,
  input         PIPELINE_RD,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         LS,
  input         SD_RB1,
  input         TEST1A,
  input         CS1,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_b0,
  input         WEN1_b1,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Full,
  output        Almost_Empty
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK2, "");
      $hold(posedge CLK2, WD_b0, "");
      $setup(WD_b1, posedge CLK2, "");
      $hold(posedge CLK2, WD_b1, "");
      $setup(WD_b2, posedge CLK2, "");
      $hold(posedge CLK2, WD_b2, "");
      $setup(WD_b3, posedge CLK2, "");
      $hold(posedge CLK2, WD_b3, "");
      $setup(WD_b4, posedge CLK2, "");
      $hold(posedge CLK2, WD_b4, "");
      $setup(WD_b5, posedge CLK2, "");
      $hold(posedge CLK2, WD_b5, "");
      $setup(WD_b6, posedge CLK2, "");
      $hold(posedge CLK2, WD_b6, "");
      $setup(WD_b7, posedge CLK2, "");
      $hold(posedge CLK2, WD_b7, "");
      $setup(WD_b8, posedge CLK2, "");
      $hold(posedge CLK2, WD_b8, "");
      $setup(WD_b9, posedge CLK2, "");
      $hold(posedge CLK2, WD_b9, "");
      $setup(WD_b10, posedge CLK2, "");
      $hold(posedge CLK2, WD_b10, "");
      $setup(WD_b11, posedge CLK2, "");
      $hold(posedge CLK2, WD_b11, "");
      $setup(WD_b12, posedge CLK2, "");
      $hold(posedge CLK2, WD_b12, "");
      $setup(WD_b13, posedge CLK2, "");
      $hold(posedge CLK2, WD_b13, "");
      $setup(WD_b14, posedge CLK2, "");
      $hold(posedge CLK2, WD_b14, "");
      $setup(WD_b15, posedge CLK2, "");
      $hold(posedge CLK2, WD_b15, "");
      $setup(WD_b16, posedge CLK2, "");
      $hold(posedge CLK2, WD_b16, "");
      $setup(WD_b17, posedge CLK2, "");
      $hold(posedge CLK2, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>POP_FLAG_b0)="";
      (CLK1*>POP_FLAG_b1)="";
      (CLK1*>POP_FLAG_b2)="";
      (CLK1*>POP_FLAG_b3)="";
      (CLK2*>PUSH_FLAG_b0)="";
      (CLK2*>PUSH_FLAG_b1)="";
      (CLK2*>PUSH_FLAG_b2)="";
      (CLK2*>PUSH_FLAG_b3)="";
      (CLK1*>RD_b0)="";
      (CLK1*>RD_b1)="";
      (CLK1*>RD_b2)="";
      (CLK1*>RD_b3)="";
      (CLK1*>RD_b4)="";
      (CLK1*>RD_b5)="";
      (CLK1*>RD_b6)="";
      (CLK1*>RD_b7)="";
      (CLK1*>RD_b8)="";
      (CLK1*>RD_b9)="";
      (CLK1*>RD_b10)="";
      (CLK1*>RD_b11)="";
      (CLK1*>RD_b12)="";
      (CLK1*>RD_b13)="";
      (CLK1*>RD_b14)="";
      (CLK1*>RD_b15)="";
      (CLK1*>RD_b16)="";
      (CLK1*>RD_b17)="";
      (CLK2*>Almost_Full)="";
      (CLK1*>Almost_Empty)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .P1_0(P1),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Full_0(Almost_Full),
      .Almost_Empty_0(Almost_Empty));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D1_PR1_WSA0_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         TEST1B,
  input         PIPELINE_RD,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         LS,
  input         SD_RB1,
  input         TEST1A,
  input         CS1,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_b0,
  input         WEN1_b1,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Full,
  output        Almost_Empty
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK2, "");
      $hold(posedge CLK2, WD_b0, "");
      $setup(WD_b1, posedge CLK2, "");
      $hold(posedge CLK2, WD_b1, "");
      $setup(WD_b2, posedge CLK2, "");
      $hold(posedge CLK2, WD_b2, "");
      $setup(WD_b3, posedge CLK2, "");
      $hold(posedge CLK2, WD_b3, "");
      $setup(WD_b4, posedge CLK2, "");
      $hold(posedge CLK2, WD_b4, "");
      $setup(WD_b5, posedge CLK2, "");
      $hold(posedge CLK2, WD_b5, "");
      $setup(WD_b6, posedge CLK2, "");
      $hold(posedge CLK2, WD_b6, "");
      $setup(WD_b7, posedge CLK2, "");
      $hold(posedge CLK2, WD_b7, "");
      $setup(WD_b8, posedge CLK2, "");
      $hold(posedge CLK2, WD_b8, "");
      $setup(WD_b9, posedge CLK2, "");
      $hold(posedge CLK2, WD_b9, "");
      $setup(WD_b10, posedge CLK2, "");
      $hold(posedge CLK2, WD_b10, "");
      $setup(WD_b11, posedge CLK2, "");
      $hold(posedge CLK2, WD_b11, "");
      $setup(WD_b12, posedge CLK2, "");
      $hold(posedge CLK2, WD_b12, "");
      $setup(WD_b13, posedge CLK2, "");
      $hold(posedge CLK2, WD_b13, "");
      $setup(WD_b14, posedge CLK2, "");
      $hold(posedge CLK2, WD_b14, "");
      $setup(WD_b15, posedge CLK2, "");
      $hold(posedge CLK2, WD_b15, "");
      $setup(WD_b16, posedge CLK2, "");
      $hold(posedge CLK2, WD_b16, "");
      $setup(WD_b17, posedge CLK2, "");
      $hold(posedge CLK2, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>POP_FLAG_b0)="";
      (CLK1*>POP_FLAG_b1)="";
      (CLK1*>POP_FLAG_b2)="";
      (CLK1*>POP_FLAG_b3)="";
      (CLK2*>PUSH_FLAG_b0)="";
      (CLK2*>PUSH_FLAG_b1)="";
      (CLK2*>PUSH_FLAG_b2)="";
      (CLK2*>PUSH_FLAG_b3)="";
      (CLK1*>RD_b0)="";
      (CLK1*>RD_b1)="";
      (CLK1*>RD_b2)="";
      (CLK1*>RD_b3)="";
      (CLK1*>RD_b4)="";
      (CLK1*>RD_b5)="";
      (CLK1*>RD_b6)="";
      (CLK1*>RD_b7)="";
      (CLK1*>RD_b8)="";
      (CLK1*>RD_b9)="";
      (CLK1*>RD_b10)="";
      (CLK1*>RD_b11)="";
      (CLK1*>RD_b12)="";
      (CLK1*>RD_b13)="";
      (CLK1*>RD_b14)="";
      (CLK1*>RD_b15)="";
      (CLK1*>RD_b16)="";
      (CLK1*>RD_b17)="";
      (CLK2*>Almost_Full)="";
      (CLK1*>Almost_Empty)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .P1_0(P1),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Full_0(Almost_Full),
      .Almost_Empty_0(Almost_Empty));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D1_PR1_WSA0_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         TEST1B,
  input         PIPELINE_RD,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         LS,
  input         SD_RB1,
  input         TEST1A,
  input         CS1,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_b0,
  input         WEN1_b1,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Full,
  output        Almost_Empty
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK2, "");
      $hold(posedge CLK2, WD_b0, "");
      $setup(WD_b1, posedge CLK2, "");
      $hold(posedge CLK2, WD_b1, "");
      $setup(WD_b2, posedge CLK2, "");
      $hold(posedge CLK2, WD_b2, "");
      $setup(WD_b3, posedge CLK2, "");
      $hold(posedge CLK2, WD_b3, "");
      $setup(WD_b4, posedge CLK2, "");
      $hold(posedge CLK2, WD_b4, "");
      $setup(WD_b5, posedge CLK2, "");
      $hold(posedge CLK2, WD_b5, "");
      $setup(WD_b6, posedge CLK2, "");
      $hold(posedge CLK2, WD_b6, "");
      $setup(WD_b7, posedge CLK2, "");
      $hold(posedge CLK2, WD_b7, "");
      $setup(WD_b8, posedge CLK2, "");
      $hold(posedge CLK2, WD_b8, "");
      $setup(WD_b9, posedge CLK2, "");
      $hold(posedge CLK2, WD_b9, "");
      $setup(WD_b10, posedge CLK2, "");
      $hold(posedge CLK2, WD_b10, "");
      $setup(WD_b11, posedge CLK2, "");
      $hold(posedge CLK2, WD_b11, "");
      $setup(WD_b12, posedge CLK2, "");
      $hold(posedge CLK2, WD_b12, "");
      $setup(WD_b13, posedge CLK2, "");
      $hold(posedge CLK2, WD_b13, "");
      $setup(WD_b14, posedge CLK2, "");
      $hold(posedge CLK2, WD_b14, "");
      $setup(WD_b15, posedge CLK2, "");
      $hold(posedge CLK2, WD_b15, "");
      $setup(WD_b16, posedge CLK2, "");
      $hold(posedge CLK2, WD_b16, "");
      $setup(WD_b17, posedge CLK2, "");
      $hold(posedge CLK2, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>POP_FLAG_b0)="";
      (CLK1*>POP_FLAG_b1)="";
      (CLK1*>POP_FLAG_b2)="";
      (CLK1*>POP_FLAG_b3)="";
      (CLK2*>PUSH_FLAG_b0)="";
      (CLK2*>PUSH_FLAG_b1)="";
      (CLK2*>PUSH_FLAG_b2)="";
      (CLK2*>PUSH_FLAG_b3)="";
      (CLK1*>RD_b0)="";
      (CLK1*>RD_b1)="";
      (CLK1*>RD_b2)="";
      (CLK1*>RD_b3)="";
      (CLK1*>RD_b4)="";
      (CLK1*>RD_b5)="";
      (CLK1*>RD_b6)="";
      (CLK1*>RD_b7)="";
      (CLK1*>RD_b8)="";
      (CLK1*>RD_b9)="";
      (CLK1*>RD_b10)="";
      (CLK1*>RD_b11)="";
      (CLK1*>RD_b12)="";
      (CLK1*>RD_b13)="";
      (CLK1*>RD_b14)="";
      (CLK1*>RD_b15)="";
      (CLK1*>RD_b16)="";
      (CLK1*>RD_b17)="";
      (CLK2*>Almost_Full)="";
      (CLK1*>Almost_Empty)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .P1_0(P1),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Full_0(Almost_Full),
      .Almost_Empty_0(Almost_Empty));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D1_PR1_WSA1_WSB0_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         TEST1B,
  input         PIPELINE_RD,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         LS,
  input         SD_RB1,
  input         TEST1A,
  input         CS1,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_b0,
  input         WEN1_b1,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Full,
  output        Almost_Empty
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK2, "");
      $hold(posedge CLK2, WD_b0, "");
      $setup(WD_b1, posedge CLK2, "");
      $hold(posedge CLK2, WD_b1, "");
      $setup(WD_b2, posedge CLK2, "");
      $hold(posedge CLK2, WD_b2, "");
      $setup(WD_b3, posedge CLK2, "");
      $hold(posedge CLK2, WD_b3, "");
      $setup(WD_b4, posedge CLK2, "");
      $hold(posedge CLK2, WD_b4, "");
      $setup(WD_b5, posedge CLK2, "");
      $hold(posedge CLK2, WD_b5, "");
      $setup(WD_b6, posedge CLK2, "");
      $hold(posedge CLK2, WD_b6, "");
      $setup(WD_b7, posedge CLK2, "");
      $hold(posedge CLK2, WD_b7, "");
      $setup(WD_b8, posedge CLK2, "");
      $hold(posedge CLK2, WD_b8, "");
      $setup(WD_b9, posedge CLK2, "");
      $hold(posedge CLK2, WD_b9, "");
      $setup(WD_b10, posedge CLK2, "");
      $hold(posedge CLK2, WD_b10, "");
      $setup(WD_b11, posedge CLK2, "");
      $hold(posedge CLK2, WD_b11, "");
      $setup(WD_b12, posedge CLK2, "");
      $hold(posedge CLK2, WD_b12, "");
      $setup(WD_b13, posedge CLK2, "");
      $hold(posedge CLK2, WD_b13, "");
      $setup(WD_b14, posedge CLK2, "");
      $hold(posedge CLK2, WD_b14, "");
      $setup(WD_b15, posedge CLK2, "");
      $hold(posedge CLK2, WD_b15, "");
      $setup(WD_b16, posedge CLK2, "");
      $hold(posedge CLK2, WD_b16, "");
      $setup(WD_b17, posedge CLK2, "");
      $hold(posedge CLK2, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>POP_FLAG_b0)="";
      (CLK1*>POP_FLAG_b1)="";
      (CLK1*>POP_FLAG_b2)="";
      (CLK1*>POP_FLAG_b3)="";
      (CLK2*>PUSH_FLAG_b0)="";
      (CLK2*>PUSH_FLAG_b1)="";
      (CLK2*>PUSH_FLAG_b2)="";
      (CLK2*>PUSH_FLAG_b3)="";
      (CLK1*>RD_b0)="";
      (CLK1*>RD_b1)="";
      (CLK1*>RD_b2)="";
      (CLK1*>RD_b3)="";
      (CLK1*>RD_b4)="";
      (CLK1*>RD_b5)="";
      (CLK1*>RD_b6)="";
      (CLK1*>RD_b7)="";
      (CLK1*>RD_b8)="";
      (CLK1*>RD_b9)="";
      (CLK1*>RD_b10)="";
      (CLK1*>RD_b11)="";
      (CLK1*>RD_b12)="";
      (CLK1*>RD_b13)="";
      (CLK1*>RD_b14)="";
      (CLK1*>RD_b15)="";
      (CLK1*>RD_b16)="";
      (CLK1*>RD_b17)="";
      (CLK2*>Almost_Full)="";
      (CLK1*>Almost_Empty)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .P1_0(P1),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Full_0(Almost_Full),
      .Almost_Empty_0(Almost_Empty));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE0_FE1_D1_PR1_WSA1_WSB1_VPR (

  input         CLK2,
  input         CLK1,

  input         DIR,
  input         DS_RB1,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         P2,
  input         FIFO_EN,
  input         CONCAT_EN,
  input         ASYNC_FLUSH,
  input         A2_b0,
  input         A2_b1,
  input         A2_b2,
  input         A2_b3,
  input         A2_b4,
  input         A2_b5,
  input         A2_b6,
  input         A2_b7,
  input         A2_b8,
  input         A2_b9,
  input         A2_b10,
  input         TEST1B,
  input         PIPELINE_RD,
  input         WD_b0,
  input         WD_b1,
  input         WD_b2,
  input         WD_b3,
  input         WD_b4,
  input         WD_b5,
  input         WD_b6,
  input         WD_b7,
  input         WD_b8,
  input         WD_b9,
  input         WD_b10,
  input         WD_b11,
  input         WD_b12,
  input         WD_b13,
  input         WD_b14,
  input         WD_b15,
  input         WD_b16,
  input         WD_b17,
  input         DS,
  input  [ 1:0] WIDTH_SELECT2,
  input         LS_RB1,
  input         CS2,
  input         LS,
  input         SD_RB1,
  input         TEST1A,
  input         CS1,
  input  [ 1:0] WIDTH_SELECT1,
  input         A1_b0,
  input         A1_b1,
  input         A1_b2,
  input         A1_b3,
  input         A1_b4,
  input         A1_b5,
  input         A1_b6,
  input         A1_b7,
  input         A1_b8,
  input         A1_b9,
  input         A1_b10,
  input         P1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_b0,
  input         WEN1_b1,
  input         RMEA,
  input         SYNC_FIFO,
  input         CLK1EN,
  input         CLK2EN,
  input         RMEB,
  input         SD,

  output        POP_FLAG_b0,
  output        POP_FLAG_b1,
  output        POP_FLAG_b2,
  output        POP_FLAG_b3,
  output        PUSH_FLAG_b0,
  output        PUSH_FLAG_b1,
  output        PUSH_FLAG_b2,
  output        PUSH_FLAG_b3,
  output        RD_b0,
  output        RD_b1,
  output        RD_b2,
  output        RD_b3,
  output        RD_b4,
  output        RD_b5,
  output        RD_b6,
  output        RD_b7,
  output        RD_b8,
  output        RD_b9,
  output        RD_b10,
  output        RD_b11,
  output        RD_b12,
  output        RD_b13,
  output        RD_b14,
  output        RD_b15,
  output        RD_b16,
  output        RD_b17,
  output        Almost_Full,
  output        Almost_Empty
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(P2, posedge CLK2, "");
      $hold(posedge CLK2, P2, "");
      $setup(WD_b0, posedge CLK2, "");
      $hold(posedge CLK2, WD_b0, "");
      $setup(WD_b1, posedge CLK2, "");
      $hold(posedge CLK2, WD_b1, "");
      $setup(WD_b2, posedge CLK2, "");
      $hold(posedge CLK2, WD_b2, "");
      $setup(WD_b3, posedge CLK2, "");
      $hold(posedge CLK2, WD_b3, "");
      $setup(WD_b4, posedge CLK2, "");
      $hold(posedge CLK2, WD_b4, "");
      $setup(WD_b5, posedge CLK2, "");
      $hold(posedge CLK2, WD_b5, "");
      $setup(WD_b6, posedge CLK2, "");
      $hold(posedge CLK2, WD_b6, "");
      $setup(WD_b7, posedge CLK2, "");
      $hold(posedge CLK2, WD_b7, "");
      $setup(WD_b8, posedge CLK2, "");
      $hold(posedge CLK2, WD_b8, "");
      $setup(WD_b9, posedge CLK2, "");
      $hold(posedge CLK2, WD_b9, "");
      $setup(WD_b10, posedge CLK2, "");
      $hold(posedge CLK2, WD_b10, "");
      $setup(WD_b11, posedge CLK2, "");
      $hold(posedge CLK2, WD_b11, "");
      $setup(WD_b12, posedge CLK2, "");
      $hold(posedge CLK2, WD_b12, "");
      $setup(WD_b13, posedge CLK2, "");
      $hold(posedge CLK2, WD_b13, "");
      $setup(WD_b14, posedge CLK2, "");
      $hold(posedge CLK2, WD_b14, "");
      $setup(WD_b15, posedge CLK2, "");
      $hold(posedge CLK2, WD_b15, "");
      $setup(WD_b16, posedge CLK2, "");
      $hold(posedge CLK2, WD_b16, "");
      $setup(WD_b17, posedge CLK2, "");
      $hold(posedge CLK2, WD_b17, "");
      $setup(P1, posedge CLK1, "");
      $hold(posedge CLK1, P1, "");
      (CLK1*>POP_FLAG_b0)="";
      (CLK1*>POP_FLAG_b1)="";
      (CLK1*>POP_FLAG_b2)="";
      (CLK1*>POP_FLAG_b3)="";
      (CLK2*>PUSH_FLAG_b0)="";
      (CLK2*>PUSH_FLAG_b1)="";
      (CLK2*>PUSH_FLAG_b2)="";
      (CLK2*>PUSH_FLAG_b3)="";
      (CLK1*>RD_b0)="";
      (CLK1*>RD_b1)="";
      (CLK1*>RD_b2)="";
      (CLK1*>RD_b3)="";
      (CLK1*>RD_b4)="";
      (CLK1*>RD_b5)="";
      (CLK1*>RD_b6)="";
      (CLK1*>RD_b7)="";
      (CLK1*>RD_b8)="";
      (CLK1*>RD_b9)="";
      (CLK1*>RD_b10)="";
      (CLK1*>RD_b11)="";
      (CLK1*>RD_b12)="";
      (CLK1*>RD_b13)="";
      (CLK1*>RD_b14)="";
      (CLK1*>RD_b15)="";
      (CLK1*>RD_b16)="";
      (CLK1*>RD_b17)="";
      (CLK2*>Almost_Full)="";
      (CLK1*>Almost_Empty)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_0(CLK2),
      .CLK1_0(CLK1),
      .DIR_0(DIR),
      .P2_0(P2),
      .FIFO_EN_0(FIFO_EN),
      .CONCAT_EN_0(CONCAT_EN),
      .ASYNC_FLUSH_0(ASYNC_FLUSH),
      .A2_0_b0(A2_b0),
      .A2_0_b1(A2_b1),
      .A2_0_b2(A2_b2),
      .A2_0_b3(A2_b3),
      .A2_0_b4(A2_b4),
      .A2_0_b5(A2_b5),
      .A2_0_b6(A2_b6),
      .A2_0_b7(A2_b7),
      .A2_0_b8(A2_b8),
      .A2_0_b9(A2_b9),
      .A2_0_b10(A2_b10),
      .PIPELINE_RD_0(PIPELINE_RD),
      .WD_0_b0(WD_b0),
      .WD_0_b1(WD_b1),
      .WD_0_b2(WD_b2),
      .WD_0_b3(WD_b3),
      .WD_0_b4(WD_b4),
      .WD_0_b5(WD_b5),
      .WD_0_b6(WD_b6),
      .WD_0_b7(WD_b7),
      .WD_0_b8(WD_b8),
      .WD_0_b9(WD_b9),
      .WD_0_b10(WD_b10),
      .WD_0_b11(WD_b11),
      .WD_0_b12(WD_b12),
      .WD_0_b13(WD_b13),
      .WD_0_b14(WD_b14),
      .WD_0_b15(WD_b15),
      .WD_0_b16(WD_b16),
      .WD_0_b17(WD_b17),
      .WIDTH_SELECT2_0(WIDTH_SELECT2),
      .CS2_0(CS2),
      .CS1_0(CS1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1),
      .A1_0_b0(A1_b0),
      .A1_0_b1(A1_b1),
      .A1_0_b2(A1_b2),
      .A1_0_b3(A1_b3),
      .A1_0_b4(A1_b4),
      .A1_0_b5(A1_b5),
      .A1_0_b6(A1_b6),
      .A1_0_b7(A1_b7),
      .A1_0_b8(A1_b8),
      .A1_0_b9(A1_b9),
      .A1_0_b10(A1_b10),
      .P1_0(P1),
      .WEN1_0_b0(WEN1_b0),
      .WEN1_0_b1(WEN1_b1),
      .SYNC_FIFO_0(SYNC_FIFO),
      .CLK1EN_0(CLK1EN),
      .CLK2EN_0(CLK2EN),
      .POP_FLAG_0_b0(POP_FLAG_b0),
      .POP_FLAG_0_b1(POP_FLAG_b1),
      .POP_FLAG_0_b2(POP_FLAG_b2),
      .POP_FLAG_0_b3(POP_FLAG_b3),
      .PUSH_FLAG_0_b0(PUSH_FLAG_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_b3),
      .RD_0_b0(RD_b0),
      .RD_0_b1(RD_b1),
      .RD_0_b2(RD_b2),
      .RD_0_b3(RD_b3),
      .RD_0_b4(RD_b4),
      .RD_0_b5(RD_b5),
      .RD_0_b6(RD_b6),
      .RD_0_b7(RD_b7),
      .RD_0_b8(RD_b8),
      .RD_0_b9(RD_b9),
      .RD_0_b10(RD_b10),
      .RD_0_b11(RD_b11),
      .RD_0_b12(RD_b12),
      .RD_0_b13(RD_b13),
      .RD_0_b14(RD_b14),
      .RD_0_b15(RD_b15),
      .RD_0_b16(RD_b16),
      .RD_0_b17(RD_b17),
      .Almost_Full_0(Almost_Full),
      .Almost_Empty_0(Almost_Empty));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR0_WSA0_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR0_WSA0_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR0_WSA0_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR0_WSA1_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR0_WSA1_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR0_WSA1_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR0_WSA2_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR0_WSA2_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR0_WSA2_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR1_WSA0_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR1_WSA0_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR1_WSA0_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR1_WSA1_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR1_WSA1_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR1_WSA1_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR1_WSA2_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR1_WSA2_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE0_PR1_WSA2_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(A1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b0, "");
      $setup(A1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b1, "");
      $setup(A1_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b2, "");
      $setup(A1_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b3, "");
      $setup(A1_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b4, "");
      $setup(A1_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b5, "");
      $setup(A1_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b6, "");
      $setup(A1_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b7, "");
      $setup(A1_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b8, "");
      $setup(A1_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b9, "");
      $setup(A1_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, A1_0_b10, "");
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(WEN1_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b0, "");
      $setup(WEN1_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WEN1_0_b1, "");
      $setup(A2_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b0, "");
      $setup(A2_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b1, "");
      $setup(A2_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b2, "");
      $setup(A2_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b3, "");
      $setup(A2_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b4, "");
      $setup(A2_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b5, "");
      $setup(A2_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b6, "");
      $setup(A2_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b7, "");
      $setup(A2_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b8, "");
      $setup(A2_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b9, "");
      $setup(A2_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, A2_0_b10, "");
      $setup(A1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b0, "");
      $setup(A1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b1, "");
      $setup(A1_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b2, "");
      $setup(A1_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b3, "");
      $setup(A1_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b4, "");
      $setup(A1_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b5, "");
      $setup(A1_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b6, "");
      $setup(A1_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b7, "");
      $setup(A1_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b8, "");
      $setup(A1_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b9, "");
      $setup(A1_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, A1_1_b10, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(WEN1_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b0, "");
      $setup(WEN1_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WEN1_1_b1, "");
      $setup(A2_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b0, "");
      $setup(A2_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b1, "");
      $setup(A2_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b2, "");
      $setup(A2_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b3, "");
      $setup(A2_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b4, "");
      $setup(A2_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b5, "");
      $setup(A2_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b6, "");
      $setup(A2_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b7, "");
      $setup(A2_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b8, "");
      $setup(A2_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b9, "");
      $setup(A2_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, A2_1_b10, "");
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR0_WSA0_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR0_WSA0_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR0_WSA0_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR0_WSA1_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR0_WSA1_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR0_WSA1_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR0_WSA2_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR0_WSA2_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR0_WSA2_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR1_WSA0_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR1_WSA0_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR1_WSA0_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR1_WSA1_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR1_WSA1_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR1_WSA1_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR1_WSA2_WSB0_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR1_WSA2_WSB1_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D0_PR1_WSA2_WSB2_VPR (

  input         CLK1_0,
  input         CLK2_0,
  input         CLK1_1,
  input         CLK2_1,

  input  [ 1:0] WIDTH_SELECT1_0,
  input         CLK1EN_0,
  input         CS1_0,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         P1_0,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         CLK2EN_0,
  input         CS2_0,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         P2_0,
  input         CONCAT_EN_0,
  input         PIPELINE_RD_0,
  input         FIFO_EN_0,
  input         DIR_0,
  input         SYNC_FIFO_0,
  input         ASYNC_FLUSH_0,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         CLK1EN_1,
  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         P1_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CLK2EN_1,
  input         CS2_1,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         P2_1,
  input         CONCAT_EN_1,
  input         PIPELINE_RD_1,
  input         FIFO_EN_1,
  input         DIR_1,
  input         SYNC_FIFO_1,
  input         ASYNC_FLUSH_1,
  input         DS,
  input         DS_RB1,
  input         LS,
  input         LS_RB1,
  input         SD,
  input         SD_RB1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         RMEA,
  input         RMEB,
  input         TEST1A,
  input         TEST1B,

  output        Almost_Full_0,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3,
  output        Almost_Empty_0,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        Almost_Full_1,
  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_1,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK1_0, "");
      $hold(posedge CLK1_0, WD_0_b17, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(WD_1_b0, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK1_1, "");
      $hold(posedge CLK1_1, WD_1_b17, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK1_0*>Almost_Full_0)="";
      (CLK1_0*>PUSH_FLAG_0_b0)="";
      (CLK1_0*>PUSH_FLAG_0_b1)="";
      (CLK1_0*>PUSH_FLAG_0_b2)="";
      (CLK1_0*>PUSH_FLAG_0_b3)="";
      (CLK2_0*>Almost_Empty_0)="";
      (CLK2_0*>POP_FLAG_0_b0)="";
      (CLK2_0*>POP_FLAG_0_b1)="";
      (CLK2_0*>POP_FLAG_0_b2)="";
      (CLK2_0*>POP_FLAG_0_b3)="";
      (CLK2_0*>RD_0_b0)="";
      (CLK2_0*>RD_0_b1)="";
      (CLK2_0*>RD_0_b2)="";
      (CLK2_0*>RD_0_b3)="";
      (CLK2_0*>RD_0_b4)="";
      (CLK2_0*>RD_0_b5)="";
      (CLK2_0*>RD_0_b6)="";
      (CLK2_0*>RD_0_b7)="";
      (CLK2_0*>RD_0_b8)="";
      (CLK2_0*>RD_0_b9)="";
      (CLK2_0*>RD_0_b10)="";
      (CLK2_0*>RD_0_b11)="";
      (CLK2_0*>RD_0_b12)="";
      (CLK2_0*>RD_0_b13)="";
      (CLK2_0*>RD_0_b14)="";
      (CLK2_0*>RD_0_b15)="";
      (CLK2_0*>RD_0_b16)="";
      (CLK2_0*>RD_0_b17)="";
      (CLK1_1*>Almost_Full_1)="";
      (CLK1_1*>PUSH_FLAG_1_b0)="";
      (CLK1_1*>PUSH_FLAG_1_b1)="";
      (CLK1_1*>PUSH_FLAG_1_b2)="";
      (CLK1_1*>PUSH_FLAG_1_b3)="";
      (CLK2_1*>Almost_Empty_1)="";
      (CLK2_1*>POP_FLAG_1_b0)="";
      (CLK2_1*>POP_FLAG_1_b1)="";
      (CLK2_1*>POP_FLAG_1_b2)="";
      (CLK2_1*>POP_FLAG_1_b3)="";
      (CLK2_1*>RD_1_b0)="";
      (CLK2_1*>RD_1_b1)="";
      (CLK2_1*>RD_1_b2)="";
      (CLK2_1*>RD_1_b3)="";
      (CLK2_1*>RD_1_b4)="";
      (CLK2_1*>RD_1_b5)="";
      (CLK2_1*>RD_1_b6)="";
      (CLK2_1*>RD_1_b7)="";
      (CLK2_1*>RD_1_b8)="";
      (CLK2_1*>RD_1_b9)="";
      (CLK2_1*>RD_1_b10)="";
      (CLK2_1*>RD_1_b11)="";
      (CLK2_1*>RD_1_b12)="";
      (CLK2_1*>RD_1_b13)="";
      (CLK2_1*>RD_1_b14)="";
      (CLK2_1*>RD_1_b15)="";
      (CLK2_1*>RD_1_b16)="";
      (CLK2_1*>RD_1_b17)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK1_0(CLK1_0),
      .CLK2_0(CLK2_0),
      .CLK1_1(CLK1_1),
      .CLK2_1(CLK2_1),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .CLK1EN_0(CLK1EN_0),
      .CS1_0(CS1_0),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .P1_0(P1_0),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .CLK2EN_0(CLK2EN_0),
      .CS2_0(CS2_0),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .P2_0(P2_0),
      .CONCAT_EN_0(CONCAT_EN_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .FIFO_EN_0(FIFO_EN_0),
      .DIR_0(DIR_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK1EN_1(CLK1EN_1),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .P1_1(P1_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CLK2EN_1(CLK2EN_1),
      .CS2_1(CS2_1),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .P2_1(P2_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .FIFO_EN_1(FIFO_EN_1),
      .DIR_1(DIR_1),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .Almost_Full_0(Almost_Full_0),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .Almost_Full_1(Almost_Full_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_1(Almost_Empty_1),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR0_WSA0_WSB0_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR0_WSA0_WSB1_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR0_WSA0_WSB2_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR0_WSA1_WSB0_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR0_WSA1_WSB1_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR0_WSA1_WSB2_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR0_WSA2_WSB0_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR0_WSA2_WSB1_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR0_WSA2_WSB2_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR1_WSA0_WSB0_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR1_WSA0_WSB1_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR1_WSA0_WSB2_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR1_WSA1_WSB0_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR1_WSA1_WSB1_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR1_WSA1_WSB2_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR1_WSA2_WSB0_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR1_WSA2_WSB1_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule

`timescale 1ns/10ps
(* blackbox *)
module RAM_CE1_FE1_D1_PR1_WSA2_WSB2_VPR (

  input         CLK2_1,
  input         CLK1_1,
  input         CLK2_0,
  input         CLK1_0,

  input         CS1_1,
  input         A1_1_b0,
  input         A1_1_b1,
  input         A1_1_b2,
  input         A1_1_b3,
  input         A1_1_b4,
  input         A1_1_b5,
  input         A1_1_b6,
  input         A1_1_b7,
  input         A1_1_b8,
  input         A1_1_b9,
  input         A1_1_b10,
  input         FIFO_EN_0,
  input         DS_RB1,
  input         CS1_0,
  input         PIPELINE_RD_0,
  input         ASYNC_FLUSH_1,
  input         DIR_1,
  input         CS2_1,
  input         CLK1EN_0,
  input  [ 1:0] WIDTH_SELECT1_0,
  input         RMB_b0,
  input         RMB_b1,
  input         RMB_b2,
  input         RMB_b3,
  input         ASYNC_FLUSH_0,
  input         SYNC_FIFO_0,
  input         SYNC_FIFO_1,
  input         RMEB,
  input         TEST1B,
  input         WD_0_b0,
  input         WD_0_b1,
  input         WD_0_b2,
  input         WD_0_b3,
  input         WD_0_b4,
  input         WD_0_b5,
  input         WD_0_b6,
  input         WD_0_b7,
  input         WD_0_b8,
  input         WD_0_b9,
  input         WD_0_b10,
  input         WD_0_b11,
  input         WD_0_b12,
  input         WD_0_b13,
  input         WD_0_b14,
  input         WD_0_b15,
  input         WD_0_b16,
  input         WD_0_b17,
  input         A2_0_b0,
  input         A2_0_b1,
  input         A2_0_b2,
  input         A2_0_b3,
  input         A2_0_b4,
  input         A2_0_b5,
  input         A2_0_b6,
  input         A2_0_b7,
  input         A2_0_b8,
  input         A2_0_b9,
  input         A2_0_b10,
  input         A1_0_b0,
  input         A1_0_b1,
  input         A1_0_b2,
  input         A1_0_b3,
  input         A1_0_b4,
  input         A1_0_b5,
  input         A1_0_b6,
  input         A1_0_b7,
  input         A1_0_b8,
  input         A1_0_b9,
  input         A1_0_b10,
  input         WEN1_1_b0,
  input         WEN1_1_b1,
  input         FIFO_EN_1,
  input         CLK2EN_0,
  input         DS,
  input         LS_RB1,
  input         CLK1EN_1,
  input  [ 1:0] WIDTH_SELECT2_0,
  input         A2_1_b0,
  input         A2_1_b1,
  input         A2_1_b2,
  input         A2_1_b3,
  input         A2_1_b4,
  input         A2_1_b5,
  input         A2_1_b6,
  input         A2_1_b7,
  input         A2_1_b8,
  input         A2_1_b9,
  input         A2_1_b10,
  input         WD_1_b0,
  input         WD_1_b1,
  input         WD_1_b2,
  input         WD_1_b3,
  input         WD_1_b4,
  input         WD_1_b5,
  input         WD_1_b6,
  input         WD_1_b7,
  input         WD_1_b8,
  input         WD_1_b9,
  input         WD_1_b10,
  input         WD_1_b11,
  input         WD_1_b12,
  input         WD_1_b13,
  input         WD_1_b14,
  input         WD_1_b15,
  input         WD_1_b16,
  input         WD_1_b17,
  input         P2_0,
  input         CS2_0,
  input         P1_1,
  input         CONCAT_EN_1,
  input         LS,
  input  [ 1:0] WIDTH_SELECT1_1,
  input         SD_RB1,
  input         TEST1A,
  input         CLK2EN_1,
  input         RMA_b0,
  input         RMA_b1,
  input         RMA_b2,
  input         RMA_b3,
  input         WEN1_0_b0,
  input         WEN1_0_b1,
  input         RMEA,
  input         DIR_0,
  input         P1_0,
  input         PIPELINE_RD_1,
  input  [ 1:0] WIDTH_SELECT2_1,
  input         CONCAT_EN_0,
  input         P2_1,
  input         SD,

  output        PUSH_FLAG_1_b0,
  output        PUSH_FLAG_1_b1,
  output        PUSH_FLAG_1_b2,
  output        PUSH_FLAG_1_b3,
  output        Almost_Empty_0,
  output        Almost_Empty_1,
  output        Almost_Full_1,
  output        RD_1_b0,
  output        RD_1_b1,
  output        RD_1_b2,
  output        RD_1_b3,
  output        RD_1_b4,
  output        RD_1_b5,
  output        RD_1_b6,
  output        RD_1_b7,
  output        RD_1_b8,
  output        RD_1_b9,
  output        RD_1_b10,
  output        RD_1_b11,
  output        RD_1_b12,
  output        RD_1_b13,
  output        RD_1_b14,
  output        RD_1_b15,
  output        RD_1_b16,
  output        RD_1_b17,
  output        Almost_Full_0,
  output        POP_FLAG_1_b0,
  output        POP_FLAG_1_b1,
  output        POP_FLAG_1_b2,
  output        POP_FLAG_1_b3,
  output        POP_FLAG_0_b0,
  output        POP_FLAG_0_b1,
  output        POP_FLAG_0_b2,
  output        POP_FLAG_0_b3,
  output        RD_0_b0,
  output        RD_0_b1,
  output        RD_0_b2,
  output        RD_0_b3,
  output        RD_0_b4,
  output        RD_0_b5,
  output        RD_0_b6,
  output        RD_0_b7,
  output        RD_0_b8,
  output        RD_0_b9,
  output        RD_0_b10,
  output        RD_0_b11,
  output        RD_0_b12,
  output        RD_0_b13,
  output        RD_0_b14,
  output        RD_0_b15,
  output        RD_0_b16,
  output        RD_0_b17,
  output        PUSH_FLAG_0_b0,
  output        PUSH_FLAG_0_b1,
  output        PUSH_FLAG_0_b2,
  output        PUSH_FLAG_0_b3
);
  parameter [18431:0] INIT = 18432'bx;

  specify
      $setup(WD_0_b0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b0, "");
      $setup(WD_0_b1, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b1, "");
      $setup(WD_0_b2, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b2, "");
      $setup(WD_0_b3, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b3, "");
      $setup(WD_0_b4, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b4, "");
      $setup(WD_0_b5, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b5, "");
      $setup(WD_0_b6, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b6, "");
      $setup(WD_0_b7, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b7, "");
      $setup(WD_0_b8, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b8, "");
      $setup(WD_0_b9, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b9, "");
      $setup(WD_0_b10, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b10, "");
      $setup(WD_0_b11, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b11, "");
      $setup(WD_0_b12, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b12, "");
      $setup(WD_0_b13, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b13, "");
      $setup(WD_0_b14, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b14, "");
      $setup(WD_0_b15, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b15, "");
      $setup(WD_0_b16, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b16, "");
      $setup(WD_0_b17, posedge CLK2_0, "");
      $hold(posedge CLK2_0, WD_0_b17, "");
      $setup(WD_1_b0, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b0, "");
      $setup(WD_1_b1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b1, "");
      $setup(WD_1_b2, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b2, "");
      $setup(WD_1_b3, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b3, "");
      $setup(WD_1_b4, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b4, "");
      $setup(WD_1_b5, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b5, "");
      $setup(WD_1_b6, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b6, "");
      $setup(WD_1_b7, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b7, "");
      $setup(WD_1_b8, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b8, "");
      $setup(WD_1_b9, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b9, "");
      $setup(WD_1_b10, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b10, "");
      $setup(WD_1_b11, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b11, "");
      $setup(WD_1_b12, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b12, "");
      $setup(WD_1_b13, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b13, "");
      $setup(WD_1_b14, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b14, "");
      $setup(WD_1_b15, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b15, "");
      $setup(WD_1_b16, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b16, "");
      $setup(WD_1_b17, posedge CLK2_1, "");
      $hold(posedge CLK2_1, WD_1_b17, "");
      $setup(P2_0, posedge CLK2_0, "");
      $hold(posedge CLK2_0, P2_0, "");
      $setup(P1_1, posedge CLK1_1, "");
      $hold(posedge CLK1_1, P1_1, "");
      $setup(P1_0, posedge CLK1_0, "");
      $hold(posedge CLK1_0, P1_0, "");
      $setup(P2_1, posedge CLK2_1, "");
      $hold(posedge CLK2_1, P2_1, "");
      (CLK2_1*>PUSH_FLAG_1_b0)="";
      (CLK2_1*>PUSH_FLAG_1_b1)="";
      (CLK2_1*>PUSH_FLAG_1_b2)="";
      (CLK2_1*>PUSH_FLAG_1_b3)="";
      (CLK1_0*>Almost_Empty_0)="";
      (CLK1_1*>Almost_Empty_1)="";
      (CLK2_1*>Almost_Full_1)="";
      (CLK1_1*>RD_1_b0)="";
      (CLK1_1*>RD_1_b1)="";
      (CLK1_1*>RD_1_b2)="";
      (CLK1_1*>RD_1_b3)="";
      (CLK1_1*>RD_1_b4)="";
      (CLK1_1*>RD_1_b5)="";
      (CLK1_1*>RD_1_b6)="";
      (CLK1_1*>RD_1_b7)="";
      (CLK1_1*>RD_1_b8)="";
      (CLK1_1*>RD_1_b9)="";
      (CLK1_1*>RD_1_b10)="";
      (CLK1_1*>RD_1_b11)="";
      (CLK1_1*>RD_1_b12)="";
      (CLK1_1*>RD_1_b13)="";
      (CLK1_1*>RD_1_b14)="";
      (CLK1_1*>RD_1_b15)="";
      (CLK1_1*>RD_1_b16)="";
      (CLK1_1*>RD_1_b17)="";
      (CLK2_0*>Almost_Full_0)="";
      (CLK1_1*>POP_FLAG_1_b0)="";
      (CLK1_1*>POP_FLAG_1_b1)="";
      (CLK1_1*>POP_FLAG_1_b2)="";
      (CLK1_1*>POP_FLAG_1_b3)="";
      (CLK1_0*>POP_FLAG_0_b0)="";
      (CLK1_0*>POP_FLAG_0_b1)="";
      (CLK1_0*>POP_FLAG_0_b2)="";
      (CLK1_0*>POP_FLAG_0_b3)="";
      (CLK1_0*>RD_0_b0)="";
      (CLK1_0*>RD_0_b1)="";
      (CLK1_0*>RD_0_b2)="";
      (CLK1_0*>RD_0_b3)="";
      (CLK1_0*>RD_0_b4)="";
      (CLK1_0*>RD_0_b5)="";
      (CLK1_0*>RD_0_b6)="";
      (CLK1_0*>RD_0_b7)="";
      (CLK1_0*>RD_0_b8)="";
      (CLK1_0*>RD_0_b9)="";
      (CLK1_0*>RD_0_b10)="";
      (CLK1_0*>RD_0_b11)="";
      (CLK1_0*>RD_0_b12)="";
      (CLK1_0*>RD_0_b13)="";
      (CLK1_0*>RD_0_b14)="";
      (CLK1_0*>RD_0_b15)="";
      (CLK1_0*>RD_0_b16)="";
      (CLK1_0*>RD_0_b17)="";
      (CLK2_0*>PUSH_FLAG_0_b0)="";
      (CLK2_0*>PUSH_FLAG_0_b1)="";
      (CLK2_0*>PUSH_FLAG_0_b2)="";
      (CLK2_0*>PUSH_FLAG_0_b3)="";
  endspecify


   ram8k_2x1_cell # (.INIT(INIT)) I1 ( 
      .CLK2_1(CLK2_1),
      .CLK1_1(CLK1_1),
      .CLK2_0(CLK2_0),
      .CLK1_0(CLK1_0),
      .CS1_1(CS1_1),
      .A1_1_b0(A1_1_b0),
      .A1_1_b1(A1_1_b1),
      .A1_1_b2(A1_1_b2),
      .A1_1_b3(A1_1_b3),
      .A1_1_b4(A1_1_b4),
      .A1_1_b5(A1_1_b5),
      .A1_1_b6(A1_1_b6),
      .A1_1_b7(A1_1_b7),
      .A1_1_b8(A1_1_b8),
      .A1_1_b9(A1_1_b9),
      .A1_1_b10(A1_1_b10),
      .FIFO_EN_0(FIFO_EN_0),
      .CS1_0(CS1_0),
      .PIPELINE_RD_0(PIPELINE_RD_0),
      .ASYNC_FLUSH_1(ASYNC_FLUSH_1),
      .DIR_1(DIR_1),
      .CS2_1(CS2_1),
      .CLK1EN_0(CLK1EN_0),
      .WIDTH_SELECT1_0(WIDTH_SELECT1_0),
      .ASYNC_FLUSH_0(ASYNC_FLUSH_0),
      .SYNC_FIFO_0(SYNC_FIFO_0),
      .SYNC_FIFO_1(SYNC_FIFO_1),
      .WD_0_b0(WD_0_b0),
      .WD_0_b1(WD_0_b1),
      .WD_0_b2(WD_0_b2),
      .WD_0_b3(WD_0_b3),
      .WD_0_b4(WD_0_b4),
      .WD_0_b5(WD_0_b5),
      .WD_0_b6(WD_0_b6),
      .WD_0_b7(WD_0_b7),
      .WD_0_b8(WD_0_b8),
      .WD_0_b9(WD_0_b9),
      .WD_0_b10(WD_0_b10),
      .WD_0_b11(WD_0_b11),
      .WD_0_b12(WD_0_b12),
      .WD_0_b13(WD_0_b13),
      .WD_0_b14(WD_0_b14),
      .WD_0_b15(WD_0_b15),
      .WD_0_b16(WD_0_b16),
      .WD_0_b17(WD_0_b17),
      .A2_0_b0(A2_0_b0),
      .A2_0_b1(A2_0_b1),
      .A2_0_b2(A2_0_b2),
      .A2_0_b3(A2_0_b3),
      .A2_0_b4(A2_0_b4),
      .A2_0_b5(A2_0_b5),
      .A2_0_b6(A2_0_b6),
      .A2_0_b7(A2_0_b7),
      .A2_0_b8(A2_0_b8),
      .A2_0_b9(A2_0_b9),
      .A2_0_b10(A2_0_b10),
      .A1_0_b0(A1_0_b0),
      .A1_0_b1(A1_0_b1),
      .A1_0_b2(A1_0_b2),
      .A1_0_b3(A1_0_b3),
      .A1_0_b4(A1_0_b4),
      .A1_0_b5(A1_0_b5),
      .A1_0_b6(A1_0_b6),
      .A1_0_b7(A1_0_b7),
      .A1_0_b8(A1_0_b8),
      .A1_0_b9(A1_0_b9),
      .A1_0_b10(A1_0_b10),
      .WEN1_1_b0(WEN1_1_b0),
      .WEN1_1_b1(WEN1_1_b1),
      .FIFO_EN_1(FIFO_EN_1),
      .CLK2EN_0(CLK2EN_0),
      .CLK1EN_1(CLK1EN_1),
      .WIDTH_SELECT2_0(WIDTH_SELECT2_0),
      .A2_1_b0(A2_1_b0),
      .A2_1_b1(A2_1_b1),
      .A2_1_b2(A2_1_b2),
      .A2_1_b3(A2_1_b3),
      .A2_1_b4(A2_1_b4),
      .A2_1_b5(A2_1_b5),
      .A2_1_b6(A2_1_b6),
      .A2_1_b7(A2_1_b7),
      .A2_1_b8(A2_1_b8),
      .A2_1_b9(A2_1_b9),
      .A2_1_b10(A2_1_b10),
      .WD_1_b0(WD_1_b0),
      .WD_1_b1(WD_1_b1),
      .WD_1_b2(WD_1_b2),
      .WD_1_b3(WD_1_b3),
      .WD_1_b4(WD_1_b4),
      .WD_1_b5(WD_1_b5),
      .WD_1_b6(WD_1_b6),
      .WD_1_b7(WD_1_b7),
      .WD_1_b8(WD_1_b8),
      .WD_1_b9(WD_1_b9),
      .WD_1_b10(WD_1_b10),
      .WD_1_b11(WD_1_b11),
      .WD_1_b12(WD_1_b12),
      .WD_1_b13(WD_1_b13),
      .WD_1_b14(WD_1_b14),
      .WD_1_b15(WD_1_b15),
      .WD_1_b16(WD_1_b16),
      .WD_1_b17(WD_1_b17),
      .P2_0(P2_0),
      .CS2_0(CS2_0),
      .P1_1(P1_1),
      .CONCAT_EN_1(CONCAT_EN_1),
      .WIDTH_SELECT1_1(WIDTH_SELECT1_1),
      .CLK2EN_1(CLK2EN_1),
      .WEN1_0_b0(WEN1_0_b0),
      .WEN1_0_b1(WEN1_0_b1),
      .DIR_0(DIR_0),
      .P1_0(P1_0),
      .PIPELINE_RD_1(PIPELINE_RD_1),
      .WIDTH_SELECT2_1(WIDTH_SELECT2_1),
      .CONCAT_EN_0(CONCAT_EN_0),
      .P2_1(P2_1),
      .PUSH_FLAG_1_b0(PUSH_FLAG_1_b0),
      .PUSH_FLAG_1_b1(PUSH_FLAG_1_b1),
      .PUSH_FLAG_1_b2(PUSH_FLAG_1_b2),
      .PUSH_FLAG_1_b3(PUSH_FLAG_1_b3),
      .Almost_Empty_0(Almost_Empty_0),
      .Almost_Empty_1(Almost_Empty_1),
      .Almost_Full_1(Almost_Full_1),
      .RD_1_b0(RD_1_b0),
      .RD_1_b1(RD_1_b1),
      .RD_1_b2(RD_1_b2),
      .RD_1_b3(RD_1_b3),
      .RD_1_b4(RD_1_b4),
      .RD_1_b5(RD_1_b5),
      .RD_1_b6(RD_1_b6),
      .RD_1_b7(RD_1_b7),
      .RD_1_b8(RD_1_b8),
      .RD_1_b9(RD_1_b9),
      .RD_1_b10(RD_1_b10),
      .RD_1_b11(RD_1_b11),
      .RD_1_b12(RD_1_b12),
      .RD_1_b13(RD_1_b13),
      .RD_1_b14(RD_1_b14),
      .RD_1_b15(RD_1_b15),
      .RD_1_b16(RD_1_b16),
      .RD_1_b17(RD_1_b17),
      .Almost_Full_0(Almost_Full_0),
      .POP_FLAG_1_b0(POP_FLAG_1_b0),
      .POP_FLAG_1_b1(POP_FLAG_1_b1),
      .POP_FLAG_1_b2(POP_FLAG_1_b2),
      .POP_FLAG_1_b3(POP_FLAG_1_b3),
      .POP_FLAG_0_b0(POP_FLAG_0_b0),
      .POP_FLAG_0_b1(POP_FLAG_0_b1),
      .POP_FLAG_0_b2(POP_FLAG_0_b2),
      .POP_FLAG_0_b3(POP_FLAG_0_b3),
      .RD_0_b0(RD_0_b0),
      .RD_0_b1(RD_0_b1),
      .RD_0_b2(RD_0_b2),
      .RD_0_b3(RD_0_b3),
      .RD_0_b4(RD_0_b4),
      .RD_0_b5(RD_0_b5),
      .RD_0_b6(RD_0_b6),
      .RD_0_b7(RD_0_b7),
      .RD_0_b8(RD_0_b8),
      .RD_0_b9(RD_0_b9),
      .RD_0_b10(RD_0_b10),
      .RD_0_b11(RD_0_b11),
      .RD_0_b12(RD_0_b12),
      .RD_0_b13(RD_0_b13),
      .RD_0_b14(RD_0_b14),
      .RD_0_b15(RD_0_b15),
      .RD_0_b16(RD_0_b16),
      .RD_0_b17(RD_0_b17),
      .PUSH_FLAG_0_b0(PUSH_FLAG_0_b0),
      .PUSH_FLAG_0_b1(PUSH_FLAG_0_b1),
      .PUSH_FLAG_0_b2(PUSH_FLAG_0_b2),
      .PUSH_FLAG_0_b3(PUSH_FLAG_0_b3));

endmodule
