------------------------------------------------------------------------
-- File : f512x8_512x8.vhd
-- Design Date: July 18,2012
-- Creation Date: Wed May 13 16:02:49 2020

-- Created By SpDE Version: SpDE 2016.2 Release
-- Author: QuickLogic Corporation,
-- Copyright (C) 1998, Customers of QuickLogic may copy and modify this
-- file for use in designing QuickLogic devices only.
-- Description : This file is autogenerated  code that describes
-- the top level design for FIFO using
-- QuickLogic's RAM block resources.
------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity f512x8_512x8 is
          port (
   DIN : in std_logic_vector (7 downto 0);
   Fifo_Push_Flush,Fifo_Pop_Flush,PUSH,POP,Clk : in std_logic;
   Clk_En,Fifo_Dir,Async_Flush : in std_logic;
   Almost_Full,Almost_Empty: out std_logic;
   PUSH_FLAG,POP_FLAG: out std_logic_vector(3 downto 0);
   DOUT : out std_logic_vector (7 downto 0));
end f512x8_512x8;

architecture arch of f512x8_512x8 is
signal GND : std_logic;
signal VCC : std_logic;
component FIFO
   generic (
             wr_depth_int:integer;
             rd_depth_int:integer;
             wr_width_int:integer;
             rd_width_int:integer;
             reg_rd_int:integer;
             sync_fifo_int:integer             );
   port( 
         DIN : in std_logic_vector (wr_width_int-1 downto 0);
         Fifo_Push_Flush,Fifo_Pop_Flush,PUSH,POP: in std_logic;
         Push_Clk,Pop_Clk: in std_logic;
         Push_Clk_En,Pop_Clk_En,Fifo_Dir,Async_Flush,Push_Clk_Sel,Pop_Clk_Sel,Async_Flush_Sel: in std_logic;
         PUSH_FLAG,POP_FLAG: out std_logic_vector(3 downto 0);
         Almost_Full,Almost_Empty: out std_logic;
         DOUT : out std_logic_vector (rd_width_int-1 downto 0));
end component ;
begin
GND <= '0';
VCC <= '1';
FIFO_INST : FIFO
Generic Map (
         wr_depth_int => 512, 
         rd_depth_int => 512,
         wr_width_int=> 8,
         rd_width_int=> 8,
         reg_rd_int => 0,
         sync_fifo_int => 1         )
Port map ( DIN=>DIN,Fifo_Push_Flush=>Fifo_Push_Flush,Fifo_Pop_Flush=>Fifo_Pop_Flush, PUSH=>PUSH,POP=>POP,
           Push_Clk=>Clk,Pop_Clk=>Clk,
           Push_Clk_En=>Clk_En,Pop_Clk_En=>Clk_En,Fifo_Dir=>Fifo_Dir,Async_Flush=>Async_Flush,Push_Clk_Sel=> GND ,Pop_Clk_Sel=> GND,Async_Flush_Sel=> GND,
           PUSH_FLAG=>PUSH_FLAG,POP_FLAG=>POP_FLAG,ALmost_Full=>Almost_Full,
           Almost_Empty=>Almost_Empty,DOUT=>DOUT);
end arch;
