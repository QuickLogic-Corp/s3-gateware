// ../../../quicklogic/pp3/primitives/vcc/vcc.sim.v {{{
(* whitebox *)
module VCC (
    output wire VCC
);

    assign VCC = 1'b1;

endmodule
// ../../../quicklogic/pp3/primitives/vcc/vcc.sim.v }}}

// ../../../quicklogic/pp3/primitives/gnd/gnd.sim.v {{{
(* whitebox *)
module GND (
    output wire GND
);

    assign GND = 1'b0;

endmodule
// ../../../quicklogic/pp3/primitives/gnd/gnd.sim.v }}}

// ../../../quicklogic/pp3/primitives/fpga_interconnect/fpga_interconnect.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
module fpga_interconnect(
		datain,
		dataout
		);
    input wire datain;
    output wire dataout;

    specify
        (datain=>dataout)=(0,0);
    endspecify

    assign dataout = datain;

endmodule
// ../../../quicklogic/pp3/primitives/fpga_interconnect/fpga_interconnect.sim.v }}}

// ../../../quicklogic/pp3/primitives/clock/clock_cell.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
module CLOCK_CELL(I_PAD, O_CLK);

    (* iopad_external_pin *)
    input  wire I_PAD;

    output wire O_CLK;
	
	specify
        (I_PAD=>O_CLK)=(0,0);
    endspecify

    assign O_CLK = I_PAD;

endmodule
// ../../../quicklogic/pp3/primitives/clock/clock_cell.sim.v }}}

// ../../../quicklogic/pp3/primitives/bidir/bidir_cell.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
module BIDIR_CELL(
    I_PAD_$inp, I_DAT, I_EN,
    O_PAD_$out, O_DAT, O_EN
);
    (* iopad_external_pin *)
    input  wire I_PAD_$inp;
    input  wire I_EN;

    input  wire O_DAT;
    input  wire O_EN;

    output wire I_DAT;

	(* iopad_external_pin *)
    output wire O_PAD_$out;
	
    specify
        (O_DAT => O_PAD_$out) = (0,0);
        (O_EN => O_PAD_$out) = (0,0);
        (I_PAD_$inp => I_DAT) = (0,0);
        (I_EN => I_DAT) = (0,0);
    endspecify
    parameter [0:0] ESEL    = 0;
    parameter [0:0] OSEL    = 0;
    parameter [0:0] FIXHOLD = 0;
    parameter [0:0] WPD     = 0;
    parameter [0:0] DS      = 0;
    assign I_DAT = (I_EN == 1'b1) ? I_PAD_$inp : 1'b0;
    assign O_PAD_$out = (O_EN == 1'b1) ? O_DAT : 1'b0;

endmodule
// ../../../quicklogic/pp3/primitives/bidir/bidir_cell.sim.v }}}

// ../../../quicklogic/pp3/primitives/sdiomux/sdiomux_cell.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
module SDIOMUX_CELL(
    I_PAD_$inp, I_DAT, I_EN,
    O_PAD_$out, O_DAT, O_EN
);
    (* iopad_external_pin *)
    input  wire I_PAD_$inp;
    input  wire I_EN;

    input  wire O_DAT;
    input  wire O_EN;

    output wire I_DAT;

    (* iopad_external_pin *)
    output wire O_PAD_$out;
	
    specify
        (O_DAT => O_PAD_$out) = (0,0);
        (O_EN => O_PAD_$out) = (0,0);
        (I_PAD_$inp => I_DAT) = (0,0);
        (I_EN => I_DAT) = (0,0);
    endspecify
    assign I_DAT = (I_EN == 1'b0) ? I_PAD_$inp : 1'b0;
    assign O_PAD_$out = (O_EN == 1'b0) ? O_DAT : 1'b0;

endmodule
// ../../../quicklogic/pp3/primitives/sdiomux/sdiomux_cell.sim.v }}}

// ../../../quicklogic/pp3/primitives/logic/t_frag.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
module T_FRAG (TBS, XAB, XSL, XA1, XA2, XB1, XB2, XZ);
    input  wire TBS;

    input  wire XAB;
    input  wire XSL;
    input  wire XA1;
    input  wire XA2;
    input  wire XB1;
    input  wire XB2;
    output wire XZ;
    
    specify
        (TBS => XZ) = (0,0);
        (XAB => XZ) = (0,0);
        (XSL => XZ) = (0,0);
        (XA1 => XZ) = (0,0);
        (XA2 => XZ) = (0,0);
        (XB1 => XZ) = (0,0);
        (XB2 => XZ) = (0,0);
    endspecify
    parameter [0:0] XAS1 = 1'b0;
    parameter [0:0] XAS2 = 1'b0;
    parameter [0:0] XBS1 = 1'b0;
    parameter [0:0] XBS2 = 1'b0;
    wire XAP1 = (XAS1) ? ~XA1 : XA1;
    wire XAP2 = (XAS2) ? ~XA2 : XA2;
    wire XBP1 = (XBS1) ? ~XB1 : XB1;
    wire XBP2 = (XBS2) ? ~XB2 : XB2;
    wire XAI = XSL ? XAP2 : XAP1;
    wire XBI = XSL ? XBP2 : XBP1;
    wire XZI = XAB ? XBI : XAI;
    assign XZ = TBS ? XZI : 1'b0;

endmodule
// ../../../quicklogic/pp3/primitives/logic/t_frag.sim.v }}}

// ../../../quicklogic/pp3/primitives/logic/b_frag.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
module B_FRAG (TBS, XAB, XSL, XA1, XA2, XB1, XB2, XZ);
    input  wire TBS;

    input  wire XAB;
    input  wire XSL;
    input  wire XA1;
    input  wire XA2;
    input  wire XB1;
    input  wire XB2;
    output wire XZ;
   
    specify
        (TBS => XZ) = (0,0);
        (XAB => XZ) = (0,0);
        (XSL => XZ) = (0,0);
        (XA1 => XZ) = (0,0);
        (XA2 => XZ) = (0,0);
        (XB1 => XZ) = (0,0);
        (XB2 => XZ) = (0,0);
    endspecify
    parameter [0:0] XAS1 = 1'b0;
    parameter [0:0] XAS2 = 1'b0;
    parameter [0:0] XBS1 = 1'b0;
    parameter [0:0] XBS2 = 1'b0;
    wire XAP1 = (XAS1) ? ~XA1 : XA1;
    wire XAP2 = (XAS2) ? ~XA2 : XA2;
    wire XBP1 = (XBS1) ? ~XB1 : XB1;
    wire XBP2 = (XBS2) ? ~XB2 : XB2;
    wire XAI = XSL ? XAP2 : XAP1;
    wire XBI = XSL ? XBP2 : XBP1;
    wire XZI = XAB ? XBI : XAI;
    assign XZ = TBS ? XZI : 1'b0;

endmodule
// ../../../quicklogic/pp3/primitives/logic/b_frag.sim.v }}}

// ../../../quicklogic/pp3/primitives/logic/q_frag.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
module Q_FRAG (QCK, QST, QRT, QEN, QZ, QD, CONST0, CONST1);
    (* clkbuf_sink *)
    input  wire QCK;
    input  wire QST;
    input  wire QRT;
    input  wire QEN;
    input  wire QD;
    (* NO_COMB *)
    input  wire CONST0;
    (* NO_COMB *)
    input  wire CONST1;
    (* CLK_TO_Q = "QCK {iopath_QCK_QZ}" *)
    output reg  QZ;
    
    specify
        (QCK => QZ) = (0,0);
        $setup(QD, posedge QCK, "");
        $hold(posedge QCK, QD, "");
        $setup(QST, posedge QCK, "");
        $hold(posedge QCK, QST, "");
        $setup(QRT, posedge QCK, "");
        $hold(posedge QCK, QRT, "");
        $setup(QEN, posedge QCK, "");
        $hold(posedge QCK, QEN, "");
        $setup(CONST0, posedge QCK, "");
        $hold(posedge QCK, CONST0, "");
        $setup(CONST1, posedge QCK, "");
        $hold(posedge QCK, CONST1, "");
    endspecify
    parameter [0:0] Z_QCKS = 1'b1;
    initial QZ <= 1'b0;

    generate if (Z_QCKS == 1'b1) begin
        always @(posedge QCK or posedge QST or posedge QRT) begin
            if (QST)
                QZ <= 1'b1;
            else if (QRT)
                QZ <= 1'b0;
            else if (QEN)
                QZ <= QD;
        end

    end else begin
        always @(negedge QCK or posedge QST or posedge QRT) begin
            if (QST)
                QZ <= 1'b1;
            else if (QRT)
                QZ <= 1'b0;
            else if (QEN)
                QZ <= QD;
        end

    end endgenerate

endmodule
// ../../../quicklogic/pp3/primitives/logic/q_frag.sim.v }}}

// ../../../quicklogic/pp3/primitives/logic/f_frag.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
module F_FRAG (F1, F2, FS, FZ);
    input  wire F1;
    input  wire F2;
    input  wire FS;

    output wire FZ;
    specify
        (F1 => FZ) = (0,0);
        (F2 => FZ) = (0,0);
        (FS => FZ) = (0,0);
    endspecify
    assign FZ = FS ? F2 : F1;

endmodule
// ../../../quicklogic/pp3/primitives/logic/f_frag.sim.v }}}

// ../../../quicklogic/pp3/primitives/logic/c_frag.sim.v {{{
(* whitebox *)
module C_FRAG (TBS, TAB, TSL, TA1, TA2, TB1, TB2, BAB, BSL, BA1, BA2, BB1, BB2, TZ, CZ);
    input  wire TBS;

    input  wire TAB;
    input  wire TSL;
    input  wire TA1;
    input  wire TA2;
    input  wire TB1;
    input  wire TB2;

    input  wire BAB;
    input  wire BSL;
    input  wire BA1;
    input  wire BA2;
    input  wire BB1;
    input  wire BB2;

    output wire TZ;

    output wire CZ;
    parameter [0:0] TAS1 = 1'b0;
    parameter [0:0] TAS2 = 1'b0;
    parameter [0:0] TBS1 = 1'b0;
    parameter [0:0] TBS2 = 1'b0;

    parameter [0:0] BAS1 = 1'b0;
    parameter [0:0] BAS2 = 1'b0;
    parameter [0:0] BBS1 = 1'b0;
    parameter [0:0] BBS2 = 1'b0;
    wire TAP1 = (TAS1) ? ~TA1 : TA1;
    wire TAP2 = (TAS2) ? ~TA2 : TA2;
    wire TBP1 = (TBS1) ? ~TB1 : TB1;
    wire TBP2 = (TBS2) ? ~TB2 : TB2;

    wire BAP1 = (BAS1) ? ~BA1 : BA1;
    wire BAP2 = (BAS2) ? ~BA2 : BA2;
    wire BBP1 = (BBS1) ? ~BB1 : BB1;
    wire BBP2 = (BBS2) ? ~BB2 : BB2;
    wire TAI = TSL ? TAP2 : TAP1;
    wire TBI = TSL ? TBP2 : TBP1;
    
    wire BAI = BSL ? BAP2 : BAP1;
    wire BBI = BSL ? BBP2 : BBP1;
    wire TZI = TAB ? TBI : TAI;
    wire BZI = BAB ? BBI : BAI;
    wire CZI = TBS ? BZI : TZI;
    assign TZ = TZI;
    assign CZ = CZI;

    specify
        (TBS => CZ) = (0,0);
        (TAB => CZ) = (0,0);
        (TSL => CZ) = (0,0);
        (TA1 => CZ) = (0,0);
        (TA2 => CZ) = (0,0);
        (TB1 => CZ) = (0,0);
        (TB2 => CZ) = (0,0);
        (BAB => CZ) = (0,0);
        (BSL => CZ) = (0,0);
        (BA1 => CZ) = (0,0);
        (BA2 => CZ) = (0,0);
        (BB1 => CZ) = (0,0);
        (BB2 => CZ) = (0,0);
        (TAB => TZ) = (0,0);
        (TSL => TZ) = (0,0);
        (TA1 => TZ) = (0,0);
        (TA2 => TZ) = (0,0);
        (TB1 => TZ) = (0,0);
        (TB2 => TZ) = (0,0);
    endspecify

endmodule
// ../../../quicklogic/pp3/primitives/logic/c_frag.sim.v }}}

// ../../../quicklogic/pp3/primitives/assp/assp.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
(* keep *)
module ASSP (
			WB_CLK,
			WBs_ACK,
			WBs_RD_DAT,
			WBs_BYTE_STB,
			WBs_CYC,
			WBs_WE,
			WBs_RD,
			WBs_STB,
			WBs_ADR,
			SDMA_Req,
			SDMA_Sreq,
			SDMA_Done,
			SDMA_Active,
			FB_msg_out,
			FB_Int_Clr,
			FB_Start,
			FB_Busy,
			WB_RST,
			Sys_PKfb_Rst,
			Sys_Clk0,
			Sys_Clk0_Rst,
			Sys_Clk1,
			Sys_Clk1_Rst,
			Sys_Pclk,
			Sys_Pclk_Rst,
			Sys_PKfb_Clk,
			FB_PKfbData,
			WBs_WR_DAT,
			FB_PKfbPush,
			FB_PKfbSOF,
			FB_PKfbEOF,
			Sensor_Int,
			FB_PKfbOverflow,
			TimeStamp,
			Sys_PSel,
			SPIm_Paddr,
			SPIm_PEnable,
			SPIm_PWrite,
			SPIm_PWdata,
			SPIm_PReady,
			SPIm_PSlvErr,
			SPIm_Prdata,
			Device_ID
			);

  input wire         WB_CLK;
  input	wire         WBs_ACK;
  input	wire  [31:0] WBs_RD_DAT;
  output wire [3:0]  WBs_BYTE_STB;
  output wire        WBs_CYC;
  output wire        WBs_WE;
  output wire        WBs_RD;
  output wire        WBs_STB;
  output wire [16:0] WBs_ADR;
  input wire  [3:0]  SDMA_Req;
  input wire  [3:0]  SDMA_Sreq;
  output wire [3:0]  SDMA_Done;
  output wire [3:0]  SDMA_Active;
  input wire  [3:0]  FB_msg_out;
  input wire  [7:0]  FB_Int_Clr;
  output wire        FB_Start;
  input wire         FB_Busy;
  output wire        WB_RST;
  output wire        Sys_PKfb_Rst;
  output wire        Sys_Clk0;
  output wire        Sys_Clk0_Rst;
  output wire        Sys_Clk1;
  output wire        Sys_Clk1_Rst;
  output wire        Sys_Pclk;
  output wire        Sys_Pclk_Rst;
  input wire         Sys_PKfb_Clk;
  input wire  [31:0] FB_PKfbData;
  output wire [31:0] WBs_WR_DAT;
  input wire  [3:0]  FB_PKfbPush;
  input wire         FB_PKfbSOF;
  input wire         FB_PKfbEOF;
  output wire [7:0]  Sensor_Int;
  
  output wire        FB_PKfbOverflow;
  
  output wire [23:0] TimeStamp;
  input wire         Sys_PSel;
  input wire  [15:0] SPIm_Paddr;
  input wire         SPIm_PEnable;
  input wire         SPIm_PWrite;
  input wire  [31:0] SPIm_PWdata;
  
  output wire        SPIm_PReady;
  
  output wire        SPIm_PSlvErr;
 
  (* DELAY_MATRIX_Sys_PSel= "{iopath_Sys_PSel_SPIm_Prdata0} {iopath_Sys_PSel_SPIm_Prdata1} {iopath_Sys_PSel_SPIm_Prdata2} {iopath_Sys_PSel_SPIm_Prdata3} {iopath_Sys_PSel_SPIm_Prdata4} {iopath_Sys_PSel_SPIm_Prdata5} {iopath_Sys_PSel_SPIm_Prdata6} {iopath_Sys_PSel_SPIm_Prdata7} {iopath_Sys_PSel_SPIm_Prdata8} {iopath_Sys_PSel_SPIm_Prdata9} {iopath_Sys_PSel_SPIm_Prdata10} {iopath_Sys_PSel_SPIm_Prdata11} {iopath_Sys_PSel_SPIm_Prdata12} {iopath_Sys_PSel_SPIm_Prdata13} {iopath_Sys_PSel_SPIm_Prdata14} {iopath_Sys_PSel_SPIm_Prdata15} {iopath_Sys_PSel_SPIm_Prdata16} {iopath_Sys_PSel_SPIm_Prdata17} {iopath_Sys_PSel_SPIm_Prdata18} {iopath_Sys_PSel_SPIm_Prdata19} {iopath_Sys_PSel_SPIm_Prdata20} {iopath_Sys_PSel_SPIm_Prdata21} {iopath_Sys_PSel_SPIm_Prdata22} {iopath_Sys_PSel_SPIm_Prdata23} {iopath_Sys_PSel_SPIm_Prdata24} {iopath_Sys_PSel_SPIm_Prdata25} {iopath_Sys_PSel_SPIm_Prdata26} {iopath_Sys_PSel_SPIm_Prdata27} {iopath_Sys_PSel_SPIm_Prdata28} {iopath_Sys_PSel_SPIm_Prdata29} {iopath_Sys_PSel_SPIm_Prdata30} {iopath_Sys_PSel_SPIm_Prdata31}" *) 
  output wire [31:0] SPIm_Prdata;
  
  input wire  [15:0] Device_ID;
  assign SPIm_Prdata = (Sys_PSel == 1'b1) ? 32'h00000000 : 32'h00000000;
  assign SPIm_PReady = (Sys_PSel == 1'b1) ? 1'b0 : 1'b0;
  assign SPIm_PSlvErr = (Sys_PSel == 1'b1) ? 1'b0 : 1'b0;
  assign FB_PKfbOverflow = (FB_PKfbPush != 4'b0000) ? 1'b0 : 1'b0;

endmodule
// ../../../quicklogic/pp3/primitives/assp/assp.sim.v }}}

// ../../../quicklogic/pp3/primitives/mult/mult.sim.v {{{
`timescale 1ns/10ps
(* whitebox *)
module MULT (
			Amult,
			Bmult,
			Valid_mult,
			Cmult,
			sel_mul_32x32
			);

	input wire  [31:0] Amult;
	input wire  [31:0] Bmult;
	input wire   [1:0] Valid_mult;
`ifndef G_SIM
`endif
	output reg  [63:0] Cmult;
	input wire         sel_mul_32x32;

`ifdef GSIM
    specify
		(Amult[0]  => Cmult[0]) = (0,0);
		(Amult[1]  => Cmult[0]) = (0,0);
		(Amult[2]  => Cmult[0]) = (0,0);
		(Amult[3]  => Cmult[0]) = (0,0);
		(Amult[4]  => Cmult[0]) = (0,0);
		(Amult[5]  => Cmult[0]) = (0,0);
		(Amult[6]  => Cmult[0]) = (0,0);
		(Amult[7]  => Cmult[0]) = (0,0);
		(Amult[8]  => Cmult[0]) = (0,0);
		(Amult[9]  => Cmult[0]) = (0,0);
		(Amult[10] => Cmult[0]) = (0,0);
		(Amult[11] => Cmult[0]) = (0,0);
		(Amult[12] => Cmult[0]) = (0,0);
		(Amult[13] => Cmult[0]) = (0,0);
		(Amult[14] => Cmult[0]) = (0,0);
		(Amult[15] => Cmult[0]) = (0,0);
		(Amult[16] => Cmult[0]) = (0,0);
		(Amult[17] => Cmult[0]) = (0,0);
		(Amult[18] => Cmult[0]) = (0,0);
		(Amult[19] => Cmult[0]) = (0,0);
		(Amult[20] => Cmult[0]) = (0,0);
		(Amult[21] => Cmult[0]) = (0,0);
		(Amult[22] => Cmult[0]) = (0,0);
		(Amult[23] => Cmult[0]) = (0,0);
		(Amult[24] => Cmult[0]) = (0,0);
		(Amult[25] => Cmult[0]) = (0,0);
		(Amult[26] => Cmult[0]) = (0,0);
		(Amult[27] => Cmult[0]) = (0,0);
		(Amult[28] => Cmult[0]) = (0,0);
		(Amult[29] => Cmult[0]) = (0,0);
		(Amult[30] => Cmult[0]) = (0,0);
		(Amult[31] => Cmult[0]) = (0,0);
		(Bmult[0]  => Cmult[0]) = (0,0);
		(Bmult[1]  => Cmult[0]) = (0,0);
		(Bmult[2]  => Cmult[0]) = (0,0);
		(Bmult[3]  => Cmult[0]) = (0,0);
		(Bmult[4]  => Cmult[0]) = (0,0);
		(Bmult[5]  => Cmult[0]) = (0,0);
		(Bmult[6]  => Cmult[0]) = (0,0);
		(Bmult[7]  => Cmult[0]) = (0,0);
		(Bmult[8]  => Cmult[0]) = (0,0);
		(Bmult[9]  => Cmult[0]) = (0,0);
		(Bmult[10] => Cmult[0]) = (0,0);
		(Bmult[11] => Cmult[0]) = (0,0);
		(Bmult[12] => Cmult[0]) = (0,0);
		(Bmult[13] => Cmult[0]) = (0,0);
		(Bmult[14] => Cmult[0]) = (0,0);
		(Bmult[15] => Cmult[0]) = (0,0);
		(Bmult[16] => Cmult[0]) = (0,0);
		(Bmult[17] => Cmult[0]) = (0,0);
		(Bmult[18] => Cmult[0]) = (0,0);
		(Bmult[19] => Cmult[0]) = (0,0);
		(Bmult[20] => Cmult[0]) = (0,0);
		(Bmult[21] => Cmult[0]) = (0,0);
		(Bmult[22] => Cmult[0]) = (0,0);
		(Bmult[23] => Cmult[0]) = (0,0);
		(Bmult[24] => Cmult[0]) = (0,0);
		(Bmult[25] => Cmult[0]) = (0,0);
		(Bmult[26] => Cmult[0]) = (0,0);
		(Bmult[27] => Cmult[0]) = (0,0);
		(Bmult[28] => Cmult[0]) = (0,0);
		(Bmult[29] => Cmult[0]) = (0,0);
		(Bmult[30] => Cmult[0]) = (0,0);
		(Bmult[31] => Cmult[0]) = (0,0);		
		(Valid_mult[0] => Cmult[0]) = (0,0);
		(Valid_mult[1] => Cmult[0]) = (0,0);
		(sel_mul_32x32 => Cmult[0]) = (0,0);
		(Amult[0]  => Cmult[1]) = (0,0);
		(Amult[1]  => Cmult[1]) = (0,0);
		(Amult[2]  => Cmult[1]) = (0,0);
		(Amult[3]  => Cmult[1]) = (0,0);
		(Amult[4]  => Cmult[1]) = (0,0);
		(Amult[5]  => Cmult[1]) = (0,0);
		(Amult[6]  => Cmult[1]) = (0,0);
		(Amult[7]  => Cmult[1]) = (0,0);
		(Amult[8]  => Cmult[1]) = (0,0);
		(Amult[9]  => Cmult[1]) = (0,0);
		(Amult[10] => Cmult[1]) = (0,0);
		(Amult[11] => Cmult[1]) = (0,0);
		(Amult[12] => Cmult[1]) = (0,0);
		(Amult[13] => Cmult[1]) = (0,0);
		(Amult[14] => Cmult[1]) = (0,0);
		(Amult[15] => Cmult[1]) = (0,0);
		(Amult[16] => Cmult[1]) = (0,0);
		(Amult[17] => Cmult[1]) = (0,0);
		(Amult[18] => Cmult[1]) = (0,0);
		(Amult[19] => Cmult[1]) = (0,0);
		(Amult[20] => Cmult[1]) = (0,0);
		(Amult[21] => Cmult[1]) = (0,0);
		(Amult[22] => Cmult[1]) = (0,0);
		(Amult[23] => Cmult[1]) = (0,0);
		(Amult[24] => Cmult[1]) = (0,0);
		(Amult[25] => Cmult[1]) = (0,0);
		(Amult[26] => Cmult[1]) = (0,0);
		(Amult[27] => Cmult[1]) = (0,0);
		(Amult[28] => Cmult[1]) = (0,0);
		(Amult[29] => Cmult[1]) = (0,0);
		(Amult[30] => Cmult[1]) = (0,0);
		(Amult[31] => Cmult[1]) = (0,0);
		(Bmult[0]  => Cmult[1]) = (0,0);
		(Bmult[1]  => Cmult[1]) = (0,0);
		(Bmult[2]  => Cmult[1]) = (0,0);
		(Bmult[3]  => Cmult[1]) = (0,0);
		(Bmult[4]  => Cmult[1]) = (0,0);
		(Bmult[5]  => Cmult[1]) = (0,0);
		(Bmult[6]  => Cmult[1]) = (0,0);
		(Bmult[7]  => Cmult[1]) = (0,0);
		(Bmult[8]  => Cmult[1]) = (0,0);
		(Bmult[9]  => Cmult[1]) = (0,0);
		(Bmult[10] => Cmult[1]) = (0,0);
		(Bmult[11] => Cmult[1]) = (0,0);
		(Bmult[12] => Cmult[1]) = (0,0);
		(Bmult[13] => Cmult[1]) = (0,0);
		(Bmult[14] => Cmult[1]) = (0,0);
		(Bmult[15] => Cmult[1]) = (0,0);
		(Bmult[16] => Cmult[1]) = (0,0);
		(Bmult[17] => Cmult[1]) = (0,0);
		(Bmult[18] => Cmult[1]) = (0,0);
		(Bmult[19] => Cmult[1]) = (0,0);
		(Bmult[20] => Cmult[1]) = (0,0);
		(Bmult[21] => Cmult[1]) = (0,0);
		(Bmult[22] => Cmult[1]) = (0,0);
		(Bmult[23] => Cmult[1]) = (0,0);
		(Bmult[24] => Cmult[1]) = (0,0);
		(Bmult[25] => Cmult[1]) = (0,0);
		(Bmult[26] => Cmult[1]) = (0,0);
		(Bmult[27] => Cmult[1]) = (0,0);
		(Bmult[28] => Cmult[1]) = (0,0);
		(Bmult[29] => Cmult[1]) = (0,0);
		(Bmult[30] => Cmult[1]) = (0,0);
		(Bmult[31] => Cmult[1]) = (0,0);		
		(Valid_mult[0] => Cmult[1]) = (0,0);
		(Valid_mult[1] => Cmult[1]) = (0,0);
		(sel_mul_32x32 => Cmult[1]) = (0,0);
		(Amult[0]  => Cmult[2]) = (0,0);
		(Amult[1]  => Cmult[2]) = (0,0);
		(Amult[2]  => Cmult[2]) = (0,0);
		(Amult[3]  => Cmult[2]) = (0,0);
		(Amult[4]  => Cmult[2]) = (0,0);
		(Amult[5]  => Cmult[2]) = (0,0);
		(Amult[6]  => Cmult[2]) = (0,0);
		(Amult[7]  => Cmult[2]) = (0,0);
		(Amult[8]  => Cmult[2]) = (0,0);
		(Amult[9]  => Cmult[2]) = (0,0);
		(Amult[10] => Cmult[2]) = (0,0);
		(Amult[11] => Cmult[2]) = (0,0);
		(Amult[12] => Cmult[2]) = (0,0);
		(Amult[13] => Cmult[2]) = (0,0);
		(Amult[14] => Cmult[2]) = (0,0);
		(Amult[15] => Cmult[2]) = (0,0);
		(Amult[16] => Cmult[2]) = (0,0);
		(Amult[17] => Cmult[2]) = (0,0);
		(Amult[18] => Cmult[2]) = (0,0);
		(Amult[19] => Cmult[2]) = (0,0);
		(Amult[20] => Cmult[2]) = (0,0);
		(Amult[21] => Cmult[2]) = (0,0);
		(Amult[22] => Cmult[2]) = (0,0);
		(Amult[23] => Cmult[2]) = (0,0);
		(Amult[24] => Cmult[2]) = (0,0);
		(Amult[25] => Cmult[2]) = (0,0);
		(Amult[26] => Cmult[2]) = (0,0);
		(Amult[27] => Cmult[2]) = (0,0);
		(Amult[28] => Cmult[2]) = (0,0);
		(Amult[29] => Cmult[2]) = (0,0);
		(Amult[30] => Cmult[2]) = (0,0);
		(Amult[31] => Cmult[2]) = (0,0);
		(Bmult[0]  => Cmult[2]) = (0,0);
		(Bmult[1]  => Cmult[2]) = (0,0);
		(Bmult[2]  => Cmult[2]) = (0,0);
		(Bmult[3]  => Cmult[2]) = (0,0);
		(Bmult[4]  => Cmult[2]) = (0,0);
		(Bmult[5]  => Cmult[2]) = (0,0);
		(Bmult[6]  => Cmult[2]) = (0,0);
		(Bmult[7]  => Cmult[2]) = (0,0);
		(Bmult[8]  => Cmult[2]) = (0,0);
		(Bmult[9]  => Cmult[2]) = (0,0);
		(Bmult[10] => Cmult[2]) = (0,0);
		(Bmult[11] => Cmult[2]) = (0,0);
		(Bmult[12] => Cmult[2]) = (0,0);
		(Bmult[13] => Cmult[2]) = (0,0);
		(Bmult[14] => Cmult[2]) = (0,0);
		(Bmult[15] => Cmult[2]) = (0,0);
		(Bmult[16] => Cmult[2]) = (0,0);
		(Bmult[17] => Cmult[2]) = (0,0);
		(Bmult[18] => Cmult[2]) = (0,0);
		(Bmult[19] => Cmult[2]) = (0,0);
		(Bmult[20] => Cmult[2]) = (0,0);
		(Bmult[21] => Cmult[2]) = (0,0);
		(Bmult[22] => Cmult[2]) = (0,0);
		(Bmult[23] => Cmult[2]) = (0,0);
		(Bmult[24] => Cmult[2]) = (0,0);
		(Bmult[25] => Cmult[2]) = (0,0);
		(Bmult[26] => Cmult[2]) = (0,0);
		(Bmult[27] => Cmult[2]) = (0,0);
		(Bmult[28] => Cmult[2]) = (0,0);
		(Bmult[29] => Cmult[2]) = (0,0);
		(Bmult[30] => Cmult[2]) = (0,0);
		(Bmult[31] => Cmult[2]) = (0,0);		
		(Valid_mult[0] => Cmult[2]) = (0,0);
		(Valid_mult[1] => Cmult[2]) = (0,0);
		(sel_mul_32x32 => Cmult[2]) = (0,0);
		(Amult[0]  => Cmult[3]) = (0,0);
		(Amult[1]  => Cmult[3]) = (0,0);
		(Amult[2]  => Cmult[3]) = (0,0);
		(Amult[3]  => Cmult[3]) = (0,0);
		(Amult[4]  => Cmult[3]) = (0,0);
		(Amult[5]  => Cmult[3]) = (0,0);
		(Amult[6]  => Cmult[3]) = (0,0);
		(Amult[7]  => Cmult[3]) = (0,0);
		(Amult[8]  => Cmult[3]) = (0,0);
		(Amult[9]  => Cmult[3]) = (0,0);
		(Amult[10] => Cmult[3]) = (0,0);
		(Amult[11] => Cmult[3]) = (0,0);
		(Amult[12] => Cmult[3]) = (0,0);
		(Amult[13] => Cmult[3]) = (0,0);
		(Amult[14] => Cmult[3]) = (0,0);
		(Amult[15] => Cmult[3]) = (0,0);
		(Amult[16] => Cmult[3]) = (0,0);
		(Amult[17] => Cmult[3]) = (0,0);
		(Amult[18] => Cmult[3]) = (0,0);
		(Amult[19] => Cmult[3]) = (0,0);
		(Amult[20] => Cmult[3]) = (0,0);
		(Amult[21] => Cmult[3]) = (0,0);
		(Amult[22] => Cmult[3]) = (0,0);
		(Amult[23] => Cmult[3]) = (0,0);
		(Amult[24] => Cmult[3]) = (0,0);
		(Amult[25] => Cmult[3]) = (0,0);
		(Amult[26] => Cmult[3]) = (0,0);
		(Amult[27] => Cmult[3]) = (0,0);
		(Amult[28] => Cmult[3]) = (0,0);
		(Amult[29] => Cmult[3]) = (0,0);
		(Amult[30] => Cmult[3]) = (0,0);
		(Amult[31] => Cmult[3]) = (0,0);
		(Bmult[0]  => Cmult[3]) = (0,0);
		(Bmult[1]  => Cmult[3]) = (0,0);
		(Bmult[2]  => Cmult[3]) = (0,0);
		(Bmult[3]  => Cmult[3]) = (0,0);
		(Bmult[4]  => Cmult[3]) = (0,0);
		(Bmult[5]  => Cmult[3]) = (0,0);
		(Bmult[6]  => Cmult[3]) = (0,0);
		(Bmult[7]  => Cmult[3]) = (0,0);
		(Bmult[8]  => Cmult[3]) = (0,0);
		(Bmult[9]  => Cmult[3]) = (0,0);
		(Bmult[10] => Cmult[3]) = (0,0);
		(Bmult[11] => Cmult[3]) = (0,0);
		(Bmult[12] => Cmult[3]) = (0,0);
		(Bmult[13] => Cmult[3]) = (0,0);
		(Bmult[14] => Cmult[3]) = (0,0);
		(Bmult[15] => Cmult[3]) = (0,0);
		(Bmult[16] => Cmult[3]) = (0,0);
		(Bmult[17] => Cmult[3]) = (0,0);
		(Bmult[18] => Cmult[3]) = (0,0);
		(Bmult[19] => Cmult[3]) = (0,0);
		(Bmult[20] => Cmult[3]) = (0,0);
		(Bmult[21] => Cmult[3]) = (0,0);
		(Bmult[22] => Cmult[3]) = (0,0);
		(Bmult[23] => Cmult[3]) = (0,0);
		(Bmult[24] => Cmult[3]) = (0,0);
		(Bmult[25] => Cmult[3]) = (0,0);
		(Bmult[26] => Cmult[3]) = (0,0);
		(Bmult[27] => Cmult[3]) = (0,0);
		(Bmult[28] => Cmult[3]) = (0,0);
		(Bmult[29] => Cmult[3]) = (0,0);
		(Bmult[30] => Cmult[3]) = (0,0);
		(Bmult[31] => Cmult[3]) = (0,0);		
		(Valid_mult[0] => Cmult[3]) = (0,0);
		(Valid_mult[1] => Cmult[3]) = (0,0);
		(sel_mul_32x32 => Cmult[3]) = (0,0);
		(Amult[0]  => Cmult[4]) = (0,0);
		(Amult[1]  => Cmult[4]) = (0,0);
		(Amult[2]  => Cmult[4]) = (0,0);
		(Amult[3]  => Cmult[4]) = (0,0);
		(Amult[4]  => Cmult[4]) = (0,0);
		(Amult[5]  => Cmult[4]) = (0,0);
		(Amult[6]  => Cmult[4]) = (0,0);
		(Amult[7]  => Cmult[4]) = (0,0);
		(Amult[8]  => Cmult[4]) = (0,0);
		(Amult[9]  => Cmult[4]) = (0,0);
		(Amult[10] => Cmult[4]) = (0,0);
		(Amult[11] => Cmult[4]) = (0,0);
		(Amult[12] => Cmult[4]) = (0,0);
		(Amult[13] => Cmult[4]) = (0,0);
		(Amult[14] => Cmult[4]) = (0,0);
		(Amult[15] => Cmult[4]) = (0,0);
		(Amult[16] => Cmult[4]) = (0,0);
		(Amult[17] => Cmult[4]) = (0,0);
		(Amult[18] => Cmult[4]) = (0,0);
		(Amult[19] => Cmult[4]) = (0,0);
		(Amult[20] => Cmult[4]) = (0,0);
		(Amult[21] => Cmult[4]) = (0,0);
		(Amult[22] => Cmult[4]) = (0,0);
		(Amult[23] => Cmult[4]) = (0,0);
		(Amult[24] => Cmult[4]) = (0,0);
		(Amult[25] => Cmult[4]) = (0,0);
		(Amult[26] => Cmult[4]) = (0,0);
		(Amult[27] => Cmult[4]) = (0,0);
		(Amult[28] => Cmult[4]) = (0,0);
		(Amult[29] => Cmult[4]) = (0,0);
		(Amult[30] => Cmult[4]) = (0,0);
		(Amult[31] => Cmult[4]) = (0,0);
		(Bmult[0]  => Cmult[4]) = (0,0);
		(Bmult[1]  => Cmult[4]) = (0,0);
		(Bmult[2]  => Cmult[4]) = (0,0);
		(Bmult[3]  => Cmult[4]) = (0,0);
		(Bmult[4]  => Cmult[4]) = (0,0);
		(Bmult[5]  => Cmult[4]) = (0,0);
		(Bmult[6]  => Cmult[4]) = (0,0);
		(Bmult[7]  => Cmult[4]) = (0,0);
		(Bmult[8]  => Cmult[4]) = (0,0);
		(Bmult[9]  => Cmult[4]) = (0,0);
		(Bmult[10] => Cmult[4]) = (0,0);
		(Bmult[11] => Cmult[4]) = (0,0);
		(Bmult[12] => Cmult[4]) = (0,0);
		(Bmult[13] => Cmult[4]) = (0,0);
		(Bmult[14] => Cmult[4]) = (0,0);
		(Bmult[15] => Cmult[4]) = (0,0);
		(Bmult[16] => Cmult[4]) = (0,0);
		(Bmult[17] => Cmult[4]) = (0,0);
		(Bmult[18] => Cmult[4]) = (0,0);
		(Bmult[19] => Cmult[4]) = (0,0);
		(Bmult[20] => Cmult[4]) = (0,0);
		(Bmult[21] => Cmult[4]) = (0,0);
		(Bmult[22] => Cmult[4]) = (0,0);
		(Bmult[23] => Cmult[4]) = (0,0);
		(Bmult[24] => Cmult[4]) = (0,0);
		(Bmult[25] => Cmult[4]) = (0,0);
		(Bmult[26] => Cmult[4]) = (0,0);
		(Bmult[27] => Cmult[4]) = (0,0);
		(Bmult[28] => Cmult[4]) = (0,0);
		(Bmult[29] => Cmult[4]) = (0,0);
		(Bmult[30] => Cmult[4]) = (0,0);
		(Bmult[31] => Cmult[4]) = (0,0);		
		(Valid_mult[0] => Cmult[4]) = (0,0);
		(Valid_mult[1] => Cmult[4]) = (0,0);
		(sel_mul_32x32 => Cmult[4]) = (0,0);
		(Amult[0]  => Cmult[5]) = (0,0);
		(Amult[1]  => Cmult[5]) = (0,0);
		(Amult[2]  => Cmult[5]) = (0,0);
		(Amult[3]  => Cmult[5]) = (0,0);
		(Amult[4]  => Cmult[5]) = (0,0);
		(Amult[5]  => Cmult[5]) = (0,0);
		(Amult[6]  => Cmult[5]) = (0,0);
		(Amult[7]  => Cmult[5]) = (0,0);
		(Amult[8]  => Cmult[5]) = (0,0);
		(Amult[9]  => Cmult[5]) = (0,0);
		(Amult[10] => Cmult[5]) = (0,0);
		(Amult[11] => Cmult[5]) = (0,0);
		(Amult[12] => Cmult[5]) = (0,0);
		(Amult[13] => Cmult[5]) = (0,0);
		(Amult[14] => Cmult[5]) = (0,0);
		(Amult[15] => Cmult[5]) = (0,0);
		(Amult[16] => Cmult[5]) = (0,0);
		(Amult[17] => Cmult[5]) = (0,0);
		(Amult[18] => Cmult[5]) = (0,0);
		(Amult[19] => Cmult[5]) = (0,0);
		(Amult[20] => Cmult[5]) = (0,0);
		(Amult[21] => Cmult[5]) = (0,0);
		(Amult[22] => Cmult[5]) = (0,0);
		(Amult[23] => Cmult[5]) = (0,0);
		(Amult[24] => Cmult[5]) = (0,0);
		(Amult[25] => Cmult[5]) = (0,0);
		(Amult[26] => Cmult[5]) = (0,0);
		(Amult[27] => Cmult[5]) = (0,0);
		(Amult[28] => Cmult[5]) = (0,0);
		(Amult[29] => Cmult[5]) = (0,0);
		(Amult[30] => Cmult[5]) = (0,0);
		(Amult[31] => Cmult[5]) = (0,0);
		(Bmult[0]  => Cmult[5]) = (0,0);
		(Bmult[1]  => Cmult[5]) = (0,0);
		(Bmult[2]  => Cmult[5]) = (0,0);
		(Bmult[3]  => Cmult[5]) = (0,0);
		(Bmult[4]  => Cmult[5]) = (0,0);
		(Bmult[5]  => Cmult[5]) = (0,0);
		(Bmult[6]  => Cmult[5]) = (0,0);
		(Bmult[7]  => Cmult[5]) = (0,0);
		(Bmult[8]  => Cmult[5]) = (0,0);
		(Bmult[9]  => Cmult[5]) = (0,0);
		(Bmult[10] => Cmult[5]) = (0,0);
		(Bmult[11] => Cmult[5]) = (0,0);
		(Bmult[12] => Cmult[5]) = (0,0);
		(Bmult[13] => Cmult[5]) = (0,0);
		(Bmult[14] => Cmult[5]) = (0,0);
		(Bmult[15] => Cmult[5]) = (0,0);
		(Bmult[16] => Cmult[5]) = (0,0);
		(Bmult[17] => Cmult[5]) = (0,0);
		(Bmult[18] => Cmult[5]) = (0,0);
		(Bmult[19] => Cmult[5]) = (0,0);
		(Bmult[20] => Cmult[5]) = (0,0);
		(Bmult[21] => Cmult[5]) = (0,0);
		(Bmult[22] => Cmult[5]) = (0,0);
		(Bmult[23] => Cmult[5]) = (0,0);
		(Bmult[24] => Cmult[5]) = (0,0);
		(Bmult[25] => Cmult[5]) = (0,0);
		(Bmult[26] => Cmult[5]) = (0,0);
		(Bmult[27] => Cmult[5]) = (0,0);
		(Bmult[28] => Cmult[5]) = (0,0);
		(Bmult[29] => Cmult[5]) = (0,0);
		(Bmult[30] => Cmult[5]) = (0,0);
		(Bmult[31] => Cmult[5]) = (0,0);		
		(Valid_mult[0] => Cmult[5]) = (0,0);
		(Valid_mult[1] => Cmult[5]) = (0,0);
		(sel_mul_32x32 => Cmult[5]) = (0,0);
		(Amult[0]  => Cmult[6]) = (0,0);
		(Amult[1]  => Cmult[6]) = (0,0);
		(Amult[2]  => Cmult[6]) = (0,0);
		(Amult[3]  => Cmult[6]) = (0,0);
		(Amult[4]  => Cmult[6]) = (0,0);
		(Amult[5]  => Cmult[6]) = (0,0);
		(Amult[6]  => Cmult[6]) = (0,0);
		(Amult[7]  => Cmult[6]) = (0,0);
		(Amult[8]  => Cmult[6]) = (0,0);
		(Amult[9]  => Cmult[6]) = (0,0);
		(Amult[10] => Cmult[6]) = (0,0);
		(Amult[11] => Cmult[6]) = (0,0);
		(Amult[12] => Cmult[6]) = (0,0);
		(Amult[13] => Cmult[6]) = (0,0);
		(Amult[14] => Cmult[6]) = (0,0);
		(Amult[15] => Cmult[6]) = (0,0);
		(Amult[16] => Cmult[6]) = (0,0);
		(Amult[17] => Cmult[6]) = (0,0);
		(Amult[18] => Cmult[6]) = (0,0);
		(Amult[19] => Cmult[6]) = (0,0);
		(Amult[20] => Cmult[6]) = (0,0);
		(Amult[21] => Cmult[6]) = (0,0);
		(Amult[22] => Cmult[6]) = (0,0);
		(Amult[23] => Cmult[6]) = (0,0);
		(Amult[24] => Cmult[6]) = (0,0);
		(Amult[25] => Cmult[6]) = (0,0);
		(Amult[26] => Cmult[6]) = (0,0);
		(Amult[27] => Cmult[6]) = (0,0);
		(Amult[28] => Cmult[6]) = (0,0);
		(Amult[29] => Cmult[6]) = (0,0);
		(Amult[30] => Cmult[6]) = (0,0);
		(Amult[31] => Cmult[6]) = (0,0);
		(Bmult[0]  => Cmult[6]) = (0,0);
		(Bmult[1]  => Cmult[6]) = (0,0);
		(Bmult[2]  => Cmult[6]) = (0,0);
		(Bmult[3]  => Cmult[6]) = (0,0);
		(Bmult[4]  => Cmult[6]) = (0,0);
		(Bmult[5]  => Cmult[6]) = (0,0);
		(Bmult[6]  => Cmult[6]) = (0,0);
		(Bmult[7]  => Cmult[6]) = (0,0);
		(Bmult[8]  => Cmult[6]) = (0,0);
		(Bmult[9]  => Cmult[6]) = (0,0);
		(Bmult[10] => Cmult[6]) = (0,0);
		(Bmult[11] => Cmult[6]) = (0,0);
		(Bmult[12] => Cmult[6]) = (0,0);
		(Bmult[13] => Cmult[6]) = (0,0);
		(Bmult[14] => Cmult[6]) = (0,0);
		(Bmult[15] => Cmult[6]) = (0,0);
		(Bmult[16] => Cmult[6]) = (0,0);
		(Bmult[17] => Cmult[6]) = (0,0);
		(Bmult[18] => Cmult[6]) = (0,0);
		(Bmult[19] => Cmult[6]) = (0,0);
		(Bmult[20] => Cmult[6]) = (0,0);
		(Bmult[21] => Cmult[6]) = (0,0);
		(Bmult[22] => Cmult[6]) = (0,0);
		(Bmult[23] => Cmult[6]) = (0,0);
		(Bmult[24] => Cmult[6]) = (0,0);
		(Bmult[25] => Cmult[6]) = (0,0);
		(Bmult[26] => Cmult[6]) = (0,0);
		(Bmult[27] => Cmult[6]) = (0,0);
		(Bmult[28] => Cmult[6]) = (0,0);
		(Bmult[29] => Cmult[6]) = (0,0);
		(Bmult[30] => Cmult[6]) = (0,0);
		(Bmult[31] => Cmult[6]) = (0,0);		
		(Valid_mult[0] => Cmult[6]) = (0,0);
		(Valid_mult[1] => Cmult[6]) = (0,0);
		(sel_mul_32x32 => Cmult[6]) = (0,0);
		(Amult[0]  => Cmult[7]) = (0,0);
		(Amult[1]  => Cmult[7]) = (0,0);
		(Amult[2]  => Cmult[7]) = (0,0);
		(Amult[3]  => Cmult[7]) = (0,0);
		(Amult[4]  => Cmult[7]) = (0,0);
		(Amult[5]  => Cmult[7]) = (0,0);
		(Amult[6]  => Cmult[7]) = (0,0);
		(Amult[7]  => Cmult[7]) = (0,0);
		(Amult[8]  => Cmult[7]) = (0,0);
		(Amult[9]  => Cmult[7]) = (0,0);
		(Amult[10] => Cmult[7]) = (0,0);
		(Amult[11] => Cmult[7]) = (0,0);
		(Amult[12] => Cmult[7]) = (0,0);
		(Amult[13] => Cmult[7]) = (0,0);
		(Amult[14] => Cmult[7]) = (0,0);
		(Amult[15] => Cmult[7]) = (0,0);
		(Amult[16] => Cmult[7]) = (0,0);
		(Amult[17] => Cmult[7]) = (0,0);
		(Amult[18] => Cmult[7]) = (0,0);
		(Amult[19] => Cmult[7]) = (0,0);
		(Amult[20] => Cmult[7]) = (0,0);
		(Amult[21] => Cmult[7]) = (0,0);
		(Amult[22] => Cmult[7]) = (0,0);
		(Amult[23] => Cmult[7]) = (0,0);
		(Amult[24] => Cmult[7]) = (0,0);
		(Amult[25] => Cmult[7]) = (0,0);
		(Amult[26] => Cmult[7]) = (0,0);
		(Amult[27] => Cmult[7]) = (0,0);
		(Amult[28] => Cmult[7]) = (0,0);
		(Amult[29] => Cmult[7]) = (0,0);
		(Amult[30] => Cmult[7]) = (0,0);
		(Amult[31] => Cmult[7]) = (0,0);
		(Bmult[0]  => Cmult[7]) = (0,0);
		(Bmult[1]  => Cmult[7]) = (0,0);
		(Bmult[2]  => Cmult[7]) = (0,0);
		(Bmult[3]  => Cmult[7]) = (0,0);
		(Bmult[4]  => Cmult[7]) = (0,0);
		(Bmult[5]  => Cmult[7]) = (0,0);
		(Bmult[6]  => Cmult[7]) = (0,0);
		(Bmult[7]  => Cmult[7]) = (0,0);
		(Bmult[8]  => Cmult[7]) = (0,0);
		(Bmult[9]  => Cmult[7]) = (0,0);
		(Bmult[10] => Cmult[7]) = (0,0);
		(Bmult[11] => Cmult[7]) = (0,0);
		(Bmult[12] => Cmult[7]) = (0,0);
		(Bmult[13] => Cmult[7]) = (0,0);
		(Bmult[14] => Cmult[7]) = (0,0);
		(Bmult[15] => Cmult[7]) = (0,0);
		(Bmult[16] => Cmult[7]) = (0,0);
		(Bmult[17] => Cmult[7]) = (0,0);
		(Bmult[18] => Cmult[7]) = (0,0);
		(Bmult[19] => Cmult[7]) = (0,0);
		(Bmult[20] => Cmult[7]) = (0,0);
		(Bmult[21] => Cmult[7]) = (0,0);
		(Bmult[22] => Cmult[7]) = (0,0);
		(Bmult[23] => Cmult[7]) = (0,0);
		(Bmult[24] => Cmult[7]) = (0,0);
		(Bmult[25] => Cmult[7]) = (0,0);
		(Bmult[26] => Cmult[7]) = (0,0);
		(Bmult[27] => Cmult[7]) = (0,0);
		(Bmult[28] => Cmult[7]) = (0,0);
		(Bmult[29] => Cmult[7]) = (0,0);
		(Bmult[30] => Cmult[7]) = (0,0);
		(Bmult[31] => Cmult[7]) = (0,0);		
		(Valid_mult[0] => Cmult[7]) = (0,0);
		(Valid_mult[1] => Cmult[7]) = (0,0);
		(sel_mul_32x32 => Cmult[7]) = (0,0);
		(Amult[0]  => Cmult[8]) = (0,0);
		(Amult[1]  => Cmult[8]) = (0,0);
		(Amult[2]  => Cmult[8]) = (0,0);
		(Amult[3]  => Cmult[8]) = (0,0);
		(Amult[4]  => Cmult[8]) = (0,0);
		(Amult[5]  => Cmult[8]) = (0,0);
		(Amult[6]  => Cmult[8]) = (0,0);
		(Amult[7]  => Cmult[8]) = (0,0);
		(Amult[8]  => Cmult[8]) = (0,0);
		(Amult[9]  => Cmult[8]) = (0,0);
		(Amult[10] => Cmult[8]) = (0,0);
		(Amult[11] => Cmult[8]) = (0,0);
		(Amult[12] => Cmult[8]) = (0,0);
		(Amult[13] => Cmult[8]) = (0,0);
		(Amult[14] => Cmult[8]) = (0,0);
		(Amult[15] => Cmult[8]) = (0,0);
		(Amult[16] => Cmult[8]) = (0,0);
		(Amult[17] => Cmult[8]) = (0,0);
		(Amult[18] => Cmult[8]) = (0,0);
		(Amult[19] => Cmult[8]) = (0,0);
		(Amult[20] => Cmult[8]) = (0,0);
		(Amult[21] => Cmult[8]) = (0,0);
		(Amult[22] => Cmult[8]) = (0,0);
		(Amult[23] => Cmult[8]) = (0,0);
		(Amult[24] => Cmult[8]) = (0,0);
		(Amult[25] => Cmult[8]) = (0,0);
		(Amult[26] => Cmult[8]) = (0,0);
		(Amult[27] => Cmult[8]) = (0,0);
		(Amult[28] => Cmult[8]) = (0,0);
		(Amult[29] => Cmult[8]) = (0,0);
		(Amult[30] => Cmult[8]) = (0,0);
		(Amult[31] => Cmult[8]) = (0,0);
		(Bmult[0]  => Cmult[8]) = (0,0);
		(Bmult[1]  => Cmult[8]) = (0,0);
		(Bmult[2]  => Cmult[8]) = (0,0);
		(Bmult[3]  => Cmult[8]) = (0,0);
		(Bmult[4]  => Cmult[8]) = (0,0);
		(Bmult[5]  => Cmult[8]) = (0,0);
		(Bmult[6]  => Cmult[8]) = (0,0);
		(Bmult[7]  => Cmult[8]) = (0,0);
		(Bmult[8]  => Cmult[8]) = (0,0);
		(Bmult[9]  => Cmult[8]) = (0,0);
		(Bmult[10] => Cmult[8]) = (0,0);
		(Bmult[11] => Cmult[8]) = (0,0);
		(Bmult[12] => Cmult[8]) = (0,0);
		(Bmult[13] => Cmult[8]) = (0,0);
		(Bmult[14] => Cmult[8]) = (0,0);
		(Bmult[15] => Cmult[8]) = (0,0);
		(Bmult[16] => Cmult[8]) = (0,0);
		(Bmult[17] => Cmult[8]) = (0,0);
		(Bmult[18] => Cmult[8]) = (0,0);
		(Bmult[19] => Cmult[8]) = (0,0);
		(Bmult[20] => Cmult[8]) = (0,0);
		(Bmult[21] => Cmult[8]) = (0,0);
		(Bmult[22] => Cmult[8]) = (0,0);
		(Bmult[23] => Cmult[8]) = (0,0);
		(Bmult[24] => Cmult[8]) = (0,0);
		(Bmult[25] => Cmult[8]) = (0,0);
		(Bmult[26] => Cmult[8]) = (0,0);
		(Bmult[27] => Cmult[8]) = (0,0);
		(Bmult[28] => Cmult[8]) = (0,0);
		(Bmult[29] => Cmult[8]) = (0,0);
		(Bmult[30] => Cmult[8]) = (0,0);
		(Bmult[31] => Cmult[8]) = (0,0);		
		(Valid_mult[0] => Cmult[8]) = (0,0);
		(Valid_mult[1] => Cmult[8]) = (0,0);
		(sel_mul_32x32 => Cmult[8]) = (0,0);	
		(Amult[0]  => Cmult[9]) = (0,0);
		(Amult[1]  => Cmult[9]) = (0,0);
		(Amult[2]  => Cmult[9]) = (0,0);
		(Amult[3]  => Cmult[9]) = (0,0);
		(Amult[4]  => Cmult[9]) = (0,0);
		(Amult[5]  => Cmult[9]) = (0,0);
		(Amult[6]  => Cmult[9]) = (0,0);
		(Amult[7]  => Cmult[9]) = (0,0);
		(Amult[8]  => Cmult[9]) = (0,0);
		(Amult[9]  => Cmult[9]) = (0,0);
		(Amult[10] => Cmult[9]) = (0,0);
		(Amult[11] => Cmult[9]) = (0,0);
		(Amult[12] => Cmult[9]) = (0,0);
		(Amult[13] => Cmult[9]) = (0,0);
		(Amult[14] => Cmult[9]) = (0,0);
		(Amult[15] => Cmult[9]) = (0,0);
		(Amult[16] => Cmult[9]) = (0,0);
		(Amult[17] => Cmult[9]) = (0,0);
		(Amult[18] => Cmult[9]) = (0,0);
		(Amult[19] => Cmult[9]) = (0,0);
		(Amult[20] => Cmult[9]) = (0,0);
		(Amult[21] => Cmult[9]) = (0,0);
		(Amult[22] => Cmult[9]) = (0,0);
		(Amult[23] => Cmult[9]) = (0,0);
		(Amult[24] => Cmult[9]) = (0,0);
		(Amult[25] => Cmult[9]) = (0,0);
		(Amult[26] => Cmult[9]) = (0,0);
		(Amult[27] => Cmult[9]) = (0,0);
		(Amult[28] => Cmult[9]) = (0,0);
		(Amult[29] => Cmult[9]) = (0,0);
		(Amult[30] => Cmult[9]) = (0,0);
		(Amult[31] => Cmult[9]) = (0,0);
		(Bmult[0]  => Cmult[9]) = (0,0);
		(Bmult[1]  => Cmult[9]) = (0,0);
		(Bmult[2]  => Cmult[9]) = (0,0);
		(Bmult[3]  => Cmult[9]) = (0,0);
		(Bmult[4]  => Cmult[9]) = (0,0);
		(Bmult[5]  => Cmult[9]) = (0,0);
		(Bmult[6]  => Cmult[9]) = (0,0);
		(Bmult[7]  => Cmult[9]) = (0,0);
		(Bmult[8]  => Cmult[9]) = (0,0);
		(Bmult[9]  => Cmult[9]) = (0,0);
		(Bmult[10] => Cmult[9]) = (0,0);
		(Bmult[11] => Cmult[9]) = (0,0);
		(Bmult[12] => Cmult[9]) = (0,0);
		(Bmult[13] => Cmult[9]) = (0,0);
		(Bmult[14] => Cmult[9]) = (0,0);
		(Bmult[15] => Cmult[9]) = (0,0);
		(Bmult[16] => Cmult[9]) = (0,0);
		(Bmult[17] => Cmult[9]) = (0,0);
		(Bmult[18] => Cmult[9]) = (0,0);
		(Bmult[19] => Cmult[9]) = (0,0);
		(Bmult[20] => Cmult[9]) = (0,0);
		(Bmult[21] => Cmult[9]) = (0,0);
		(Bmult[22] => Cmult[9]) = (0,0);
		(Bmult[23] => Cmult[9]) = (0,0);
		(Bmult[24] => Cmult[9]) = (0,0);
		(Bmult[25] => Cmult[9]) = (0,0);
		(Bmult[26] => Cmult[9]) = (0,0);
		(Bmult[27] => Cmult[9]) = (0,0);
		(Bmult[28] => Cmult[9]) = (0,0);
		(Bmult[29] => Cmult[9]) = (0,0);
		(Bmult[30] => Cmult[9]) = (0,0);
		(Bmult[31] => Cmult[9]) = (0,0);		
		(Valid_mult[0] => Cmult[9]) = (0,0);
		(Valid_mult[1] => Cmult[9]) = (0,0);
		(sel_mul_32x32 => Cmult[9]) = (0,0);	
		(Amult[0]  => Cmult[10]) = (0,0);
		(Amult[1]  => Cmult[10]) = (0,0);
		(Amult[2]  => Cmult[10]) = (0,0);
		(Amult[3]  => Cmult[10]) = (0,0);
		(Amult[4]  => Cmult[10]) = (0,0);
		(Amult[5]  => Cmult[10]) = (0,0);
		(Amult[6]  => Cmult[10]) = (0,0);
		(Amult[7]  => Cmult[10]) = (0,0);
		(Amult[8]  => Cmult[10]) = (0,0);
		(Amult[9]  => Cmult[10]) = (0,0);
		(Amult[10] => Cmult[10]) = (0,0);
		(Amult[11] => Cmult[10]) = (0,0);
		(Amult[12] => Cmult[10]) = (0,0);
		(Amult[13] => Cmult[10]) = (0,0);
		(Amult[14] => Cmult[10]) = (0,0);
		(Amult[15] => Cmult[10]) = (0,0);
		(Amult[16] => Cmult[10]) = (0,0);
		(Amult[17] => Cmult[10]) = (0,0);
		(Amult[18] => Cmult[10]) = (0,0);
		(Amult[19] => Cmult[10]) = (0,0);
		(Amult[20] => Cmult[10]) = (0,0);
		(Amult[21] => Cmult[10]) = (0,0);
		(Amult[22] => Cmult[10]) = (0,0);
		(Amult[23] => Cmult[10]) = (0,0);
		(Amult[24] => Cmult[10]) = (0,0);
		(Amult[25] => Cmult[10]) = (0,0);
		(Amult[26] => Cmult[10]) = (0,0);
		(Amult[27] => Cmult[10]) = (0,0);
		(Amult[28] => Cmult[10]) = (0,0);
		(Amult[29] => Cmult[10]) = (0,0);
		(Amult[30] => Cmult[10]) = (0,0);
		(Amult[31] => Cmult[10]) = (0,0);
		(Bmult[0]  => Cmult[10]) = (0,0);
		(Bmult[1]  => Cmult[10]) = (0,0);
		(Bmult[2]  => Cmult[10]) = (0,0);
		(Bmult[3]  => Cmult[10]) = (0,0);
		(Bmult[4]  => Cmult[10]) = (0,0);
		(Bmult[5]  => Cmult[10]) = (0,0);
		(Bmult[6]  => Cmult[10]) = (0,0);
		(Bmult[7]  => Cmult[10]) = (0,0);
		(Bmult[8]  => Cmult[10]) = (0,0);
		(Bmult[9]  => Cmult[10]) = (0,0);
		(Bmult[10] => Cmult[10]) = (0,0);
		(Bmult[11] => Cmult[10]) = (0,0);
		(Bmult[12] => Cmult[10]) = (0,0);
		(Bmult[13] => Cmult[10]) = (0,0);
		(Bmult[14] => Cmult[10]) = (0,0);
		(Bmult[15] => Cmult[10]) = (0,0);
		(Bmult[16] => Cmult[10]) = (0,0);
		(Bmult[17] => Cmult[10]) = (0,0);
		(Bmult[18] => Cmult[10]) = (0,0);
		(Bmult[19] => Cmult[10]) = (0,0);
		(Bmult[20] => Cmult[10]) = (0,0);
		(Bmult[21] => Cmult[10]) = (0,0);
		(Bmult[22] => Cmult[10]) = (0,0);
		(Bmult[23] => Cmult[10]) = (0,0);
		(Bmult[24] => Cmult[10]) = (0,0);
		(Bmult[25] => Cmult[10]) = (0,0);
		(Bmult[26] => Cmult[10]) = (0,0);
		(Bmult[27] => Cmult[10]) = (0,0);
		(Bmult[28] => Cmult[10]) = (0,0);
		(Bmult[29] => Cmult[10]) = (0,0);
		(Bmult[30] => Cmult[10]) = (0,0);
		(Bmult[31] => Cmult[10]) = (0,0);		
		(Valid_mult[0] => Cmult[10]) = (0,0);
		(Valid_mult[1] => Cmult[10]) = (0,0);
		(sel_mul_32x32 => Cmult[10]) = (0,0);
		(Amult[0]  => Cmult[11]) = (0,0);
		(Amult[1]  => Cmult[11]) = (0,0);
		(Amult[2]  => Cmult[11]) = (0,0);
		(Amult[3]  => Cmult[11]) = (0,0);
		(Amult[4]  => Cmult[11]) = (0,0);
		(Amult[5]  => Cmult[11]) = (0,0);
		(Amult[6]  => Cmult[11]) = (0,0);
		(Amult[7]  => Cmult[11]) = (0,0);
		(Amult[8]  => Cmult[11]) = (0,0);
		(Amult[9]  => Cmult[11]) = (0,0);
		(Amult[10] => Cmult[11]) = (0,0);
		(Amult[11] => Cmult[11]) = (0,0);
		(Amult[12] => Cmult[11]) = (0,0);
		(Amult[13] => Cmult[11]) = (0,0);
		(Amult[14] => Cmult[11]) = (0,0);
		(Amult[15] => Cmult[11]) = (0,0);
		(Amult[16] => Cmult[11]) = (0,0);
		(Amult[17] => Cmult[11]) = (0,0);
		(Amult[18] => Cmult[11]) = (0,0);
		(Amult[19] => Cmult[11]) = (0,0);
		(Amult[20] => Cmult[11]) = (0,0);
		(Amult[21] => Cmult[11]) = (0,0);
		(Amult[22] => Cmult[11]) = (0,0);
		(Amult[23] => Cmult[11]) = (0,0);
		(Amult[24] => Cmult[11]) = (0,0);
		(Amult[25] => Cmult[11]) = (0,0);
		(Amult[26] => Cmult[11]) = (0,0);
		(Amult[27] => Cmult[11]) = (0,0);
		(Amult[28] => Cmult[11]) = (0,0);
		(Amult[29] => Cmult[11]) = (0,0);
		(Amult[30] => Cmult[11]) = (0,0);
		(Amult[31] => Cmult[11]) = (0,0);
		(Bmult[0]  => Cmult[11]) = (0,0);
		(Bmult[1]  => Cmult[11]) = (0,0);
		(Bmult[2]  => Cmult[11]) = (0,0);
		(Bmult[3]  => Cmult[11]) = (0,0);
		(Bmult[4]  => Cmult[11]) = (0,0);
		(Bmult[5]  => Cmult[11]) = (0,0);
		(Bmult[6]  => Cmult[11]) = (0,0);
		(Bmult[7]  => Cmult[11]) = (0,0);
		(Bmult[8]  => Cmult[11]) = (0,0);
		(Bmult[9]  => Cmult[11]) = (0,0);
		(Bmult[10] => Cmult[11]) = (0,0);
		(Bmult[11] => Cmult[11]) = (0,0);
		(Bmult[12] => Cmult[11]) = (0,0);
		(Bmult[13] => Cmult[11]) = (0,0);
		(Bmult[14] => Cmult[11]) = (0,0);
		(Bmult[15] => Cmult[11]) = (0,0);
		(Bmult[16] => Cmult[11]) = (0,0);
		(Bmult[17] => Cmult[11]) = (0,0);
		(Bmult[18] => Cmult[11]) = (0,0);
		(Bmult[19] => Cmult[11]) = (0,0);
		(Bmult[20] => Cmult[11]) = (0,0);
		(Bmult[21] => Cmult[11]) = (0,0);
		(Bmult[22] => Cmult[11]) = (0,0);
		(Bmult[23] => Cmult[11]) = (0,0);
		(Bmult[24] => Cmult[11]) = (0,0);
		(Bmult[25] => Cmult[11]) = (0,0);
		(Bmult[26] => Cmult[11]) = (0,0);
		(Bmult[27] => Cmult[11]) = (0,0);
		(Bmult[28] => Cmult[11]) = (0,0);
		(Bmult[29] => Cmult[11]) = (0,0);
		(Bmult[30] => Cmult[11]) = (0,0);
		(Bmult[31] => Cmult[11]) = (0,0);		
		(Valid_mult[0] => Cmult[11]) = (0,0);
		(Valid_mult[1] => Cmult[11]) = (0,0);
		(sel_mul_32x32 => Cmult[11]) = (0,0);
		(Amult[0]  => Cmult[12]) = (0,0);
		(Amult[1]  => Cmult[12]) = (0,0);
		(Amult[2]  => Cmult[12]) = (0,0);
		(Amult[3]  => Cmult[12]) = (0,0);
		(Amult[4]  => Cmult[12]) = (0,0);
		(Amult[5]  => Cmult[12]) = (0,0);
		(Amult[6]  => Cmult[12]) = (0,0);
		(Amult[7]  => Cmult[12]) = (0,0);
		(Amult[8]  => Cmult[12]) = (0,0);
		(Amult[9]  => Cmult[12]) = (0,0);
		(Amult[10] => Cmult[12]) = (0,0);
		(Amult[11] => Cmult[12]) = (0,0);
		(Amult[12] => Cmult[12]) = (0,0);
		(Amult[13] => Cmult[12]) = (0,0);
		(Amult[14] => Cmult[12]) = (0,0);
		(Amult[15] => Cmult[12]) = (0,0);
		(Amult[16] => Cmult[12]) = (0,0);
		(Amult[17] => Cmult[12]) = (0,0);
		(Amult[18] => Cmult[12]) = (0,0);
		(Amult[19] => Cmult[12]) = (0,0);
		(Amult[20] => Cmult[12]) = (0,0);
		(Amult[21] => Cmult[12]) = (0,0);
		(Amult[22] => Cmult[12]) = (0,0);
		(Amult[23] => Cmult[12]) = (0,0);
		(Amult[24] => Cmult[12]) = (0,0);
		(Amult[25] => Cmult[12]) = (0,0);
		(Amult[26] => Cmult[12]) = (0,0);
		(Amult[27] => Cmult[12]) = (0,0);
		(Amult[28] => Cmult[12]) = (0,0);
		(Amult[29] => Cmult[12]) = (0,0);
		(Amult[30] => Cmult[12]) = (0,0);
		(Amult[31] => Cmult[12]) = (0,0);
		(Bmult[0]  => Cmult[12]) = (0,0);
		(Bmult[1]  => Cmult[12]) = (0,0);
		(Bmult[2]  => Cmult[12]) = (0,0);
		(Bmult[3]  => Cmult[12]) = (0,0);
		(Bmult[4]  => Cmult[12]) = (0,0);
		(Bmult[5]  => Cmult[12]) = (0,0);
		(Bmult[6]  => Cmult[12]) = (0,0);
		(Bmult[7]  => Cmult[12]) = (0,0);
		(Bmult[8]  => Cmult[12]) = (0,0);
		(Bmult[9]  => Cmult[12]) = (0,0);
		(Bmult[10] => Cmult[12]) = (0,0);
		(Bmult[11] => Cmult[12]) = (0,0);
		(Bmult[12] => Cmult[12]) = (0,0);
		(Bmult[13] => Cmult[12]) = (0,0);
		(Bmult[14] => Cmult[12]) = (0,0);
		(Bmult[15] => Cmult[12]) = (0,0);
		(Bmult[16] => Cmult[12]) = (0,0);
		(Bmult[17] => Cmult[12]) = (0,0);
		(Bmult[18] => Cmult[12]) = (0,0);
		(Bmult[19] => Cmult[12]) = (0,0);
		(Bmult[20] => Cmult[12]) = (0,0);
		(Bmult[21] => Cmult[12]) = (0,0);
		(Bmult[22] => Cmult[12]) = (0,0);
		(Bmult[23] => Cmult[12]) = (0,0);
		(Bmult[24] => Cmult[12]) = (0,0);
		(Bmult[25] => Cmult[12]) = (0,0);
		(Bmult[26] => Cmult[12]) = (0,0);
		(Bmult[27] => Cmult[12]) = (0,0);
		(Bmult[28] => Cmult[12]) = (0,0);
		(Bmult[29] => Cmult[12]) = (0,0);
		(Bmult[30] => Cmult[12]) = (0,0);
		(Bmult[31] => Cmult[12]) = (0,0);		
		(Valid_mult[0] => Cmult[12]) = (0,0);
		(Valid_mult[1] => Cmult[12]) = (0,0);
		(sel_mul_32x32 => Cmult[12]) = (0,0);
		(Amult[0]  => Cmult[13]) = (0,0);
		(Amult[1]  => Cmult[13]) = (0,0);
		(Amult[2]  => Cmult[13]) = (0,0);
		(Amult[3]  => Cmult[13]) = (0,0);
		(Amult[4]  => Cmult[13]) = (0,0);
		(Amult[5]  => Cmult[13]) = (0,0);
		(Amult[6]  => Cmult[13]) = (0,0);
		(Amult[7]  => Cmult[13]) = (0,0);
		(Amult[8]  => Cmult[13]) = (0,0);
		(Amult[9]  => Cmult[13]) = (0,0);
		(Amult[10] => Cmult[13]) = (0,0);
		(Amult[11] => Cmult[13]) = (0,0);
		(Amult[12] => Cmult[13]) = (0,0);
		(Amult[13] => Cmult[13]) = (0,0);
		(Amult[14] => Cmult[13]) = (0,0);
		(Amult[15] => Cmult[13]) = (0,0);
		(Amult[16] => Cmult[13]) = (0,0);
		(Amult[17] => Cmult[13]) = (0,0);
		(Amult[18] => Cmult[13]) = (0,0);
		(Amult[19] => Cmult[13]) = (0,0);
		(Amult[20] => Cmult[13]) = (0,0);
		(Amult[21] => Cmult[13]) = (0,0);
		(Amult[22] => Cmult[13]) = (0,0);
		(Amult[23] => Cmult[13]) = (0,0);
		(Amult[24] => Cmult[13]) = (0,0);
		(Amult[25] => Cmult[13]) = (0,0);
		(Amult[26] => Cmult[13]) = (0,0);
		(Amult[27] => Cmult[13]) = (0,0);
		(Amult[28] => Cmult[13]) = (0,0);
		(Amult[29] => Cmult[13]) = (0,0);
		(Amult[30] => Cmult[13]) = (0,0);
		(Amult[31] => Cmult[13]) = (0,0);
		(Bmult[0]  => Cmult[13]) = (0,0);
		(Bmult[1]  => Cmult[13]) = (0,0);
		(Bmult[2]  => Cmult[13]) = (0,0);
		(Bmult[3]  => Cmult[13]) = (0,0);
		(Bmult[4]  => Cmult[13]) = (0,0);
		(Bmult[5]  => Cmult[13]) = (0,0);
		(Bmult[6]  => Cmult[13]) = (0,0);
		(Bmult[7]  => Cmult[13]) = (0,0);
		(Bmult[8]  => Cmult[13]) = (0,0);
		(Bmult[9]  => Cmult[13]) = (0,0);
		(Bmult[10] => Cmult[13]) = (0,0);
		(Bmult[11] => Cmult[13]) = (0,0);
		(Bmult[12] => Cmult[13]) = (0,0);
		(Bmult[13] => Cmult[13]) = (0,0);
		(Bmult[14] => Cmult[13]) = (0,0);
		(Bmult[15] => Cmult[13]) = (0,0);
		(Bmult[16] => Cmult[13]) = (0,0);
		(Bmult[17] => Cmult[13]) = (0,0);
		(Bmult[18] => Cmult[13]) = (0,0);
		(Bmult[19] => Cmult[13]) = (0,0);
		(Bmult[20] => Cmult[13]) = (0,0);
		(Bmult[21] => Cmult[13]) = (0,0);
		(Bmult[22] => Cmult[13]) = (0,0);
		(Bmult[23] => Cmult[13]) = (0,0);
		(Bmult[24] => Cmult[13]) = (0,0);
		(Bmult[25] => Cmult[13]) = (0,0);
		(Bmult[26] => Cmult[13]) = (0,0);
		(Bmult[27] => Cmult[13]) = (0,0);
		(Bmult[28] => Cmult[13]) = (0,0);
		(Bmult[29] => Cmult[13]) = (0,0);
		(Bmult[30] => Cmult[13]) = (0,0);
		(Bmult[31] => Cmult[13]) = (0,0);		
		(Valid_mult[0] => Cmult[13]) = (0,0);
		(Valid_mult[1] => Cmult[13]) = (0,0);
		(sel_mul_32x32 => Cmult[13]) = (0,0);
		(Amult[0]  => Cmult[14]) = (0,0);
		(Amult[1]  => Cmult[14]) = (0,0);
		(Amult[2]  => Cmult[14]) = (0,0);
		(Amult[3]  => Cmult[14]) = (0,0);
		(Amult[4]  => Cmult[14]) = (0,0);
		(Amult[5]  => Cmult[14]) = (0,0);
		(Amult[6]  => Cmult[14]) = (0,0);
		(Amult[7]  => Cmult[14]) = (0,0);
		(Amult[8]  => Cmult[14]) = (0,0);
		(Amult[9]  => Cmult[14]) = (0,0);
		(Amult[10] => Cmult[14]) = (0,0);
		(Amult[11] => Cmult[14]) = (0,0);
		(Amult[12] => Cmult[14]) = (0,0);
		(Amult[13] => Cmult[14]) = (0,0);
		(Amult[14] => Cmult[14]) = (0,0);
		(Amult[15] => Cmult[14]) = (0,0);
		(Amult[16] => Cmult[14]) = (0,0);
		(Amult[17] => Cmult[14]) = (0,0);
		(Amult[18] => Cmult[14]) = (0,0);
		(Amult[19] => Cmult[14]) = (0,0);
		(Amult[20] => Cmult[14]) = (0,0);
		(Amult[21] => Cmult[14]) = (0,0);
		(Amult[22] => Cmult[14]) = (0,0);
		(Amult[23] => Cmult[14]) = (0,0);
		(Amult[24] => Cmult[14]) = (0,0);
		(Amult[25] => Cmult[14]) = (0,0);
		(Amult[26] => Cmult[14]) = (0,0);
		(Amult[27] => Cmult[14]) = (0,0);
		(Amult[28] => Cmult[14]) = (0,0);
		(Amult[29] => Cmult[14]) = (0,0);
		(Amult[30] => Cmult[14]) = (0,0);
		(Amult[31] => Cmult[14]) = (0,0);
		(Bmult[0]  => Cmult[14]) = (0,0);
		(Bmult[1]  => Cmult[14]) = (0,0);
		(Bmult[2]  => Cmult[14]) = (0,0);
		(Bmult[3]  => Cmult[14]) = (0,0);
		(Bmult[4]  => Cmult[14]) = (0,0);
		(Bmult[5]  => Cmult[14]) = (0,0);
		(Bmult[6]  => Cmult[14]) = (0,0);
		(Bmult[7]  => Cmult[14]) = (0,0);
		(Bmult[8]  => Cmult[14]) = (0,0);
		(Bmult[9]  => Cmult[14]) = (0,0);
		(Bmult[10] => Cmult[14]) = (0,0);
		(Bmult[11] => Cmult[14]) = (0,0);
		(Bmult[12] => Cmult[14]) = (0,0);
		(Bmult[13] => Cmult[14]) = (0,0);
		(Bmult[14] => Cmult[14]) = (0,0);
		(Bmult[15] => Cmult[14]) = (0,0);
		(Bmult[16] => Cmult[14]) = (0,0);
		(Bmult[17] => Cmult[14]) = (0,0);
		(Bmult[18] => Cmult[14]) = (0,0);
		(Bmult[19] => Cmult[14]) = (0,0);
		(Bmult[20] => Cmult[14]) = (0,0);
		(Bmult[21] => Cmult[14]) = (0,0);
		(Bmult[22] => Cmult[14]) = (0,0);
		(Bmult[23] => Cmult[14]) = (0,0);
		(Bmult[24] => Cmult[14]) = (0,0);
		(Bmult[25] => Cmult[14]) = (0,0);
		(Bmult[26] => Cmult[14]) = (0,0);
		(Bmult[27] => Cmult[14]) = (0,0);
		(Bmult[28] => Cmult[14]) = (0,0);
		(Bmult[29] => Cmult[14]) = (0,0);
		(Bmult[30] => Cmult[14]) = (0,0);
		(Bmult[31] => Cmult[14]) = (0,0);		
		(Valid_mult[0] => Cmult[14]) = (0,0);
		(Valid_mult[1] => Cmult[14]) = (0,0);
		(sel_mul_32x32 => Cmult[14]) = (0,0);
		(Amult[0]  => Cmult[15]) = (0,0);
		(Amult[1]  => Cmult[15]) = (0,0);
		(Amult[2]  => Cmult[15]) = (0,0);
		(Amult[3]  => Cmult[15]) = (0,0);
		(Amult[4]  => Cmult[15]) = (0,0);
		(Amult[5]  => Cmult[15]) = (0,0);
		(Amult[6]  => Cmult[15]) = (0,0);
		(Amult[7]  => Cmult[15]) = (0,0);
		(Amult[8]  => Cmult[15]) = (0,0);
		(Amult[9]  => Cmult[15]) = (0,0);
		(Amult[10] => Cmult[15]) = (0,0);
		(Amult[11] => Cmult[15]) = (0,0);
		(Amult[12] => Cmult[15]) = (0,0);
		(Amult[13] => Cmult[15]) = (0,0);
		(Amult[14] => Cmult[15]) = (0,0);
		(Amult[15] => Cmult[15]) = (0,0);
		(Amult[16] => Cmult[15]) = (0,0);
		(Amult[17] => Cmult[15]) = (0,0);
		(Amult[18] => Cmult[15]) = (0,0);
		(Amult[19] => Cmult[15]) = (0,0);
		(Amult[20] => Cmult[15]) = (0,0);
		(Amult[21] => Cmult[15]) = (0,0);
		(Amult[22] => Cmult[15]) = (0,0);
		(Amult[23] => Cmult[15]) = (0,0);
		(Amult[24] => Cmult[15]) = (0,0);
		(Amult[25] => Cmult[15]) = (0,0);
		(Amult[26] => Cmult[15]) = (0,0);
		(Amult[27] => Cmult[15]) = (0,0);
		(Amult[28] => Cmult[15]) = (0,0);
		(Amult[29] => Cmult[15]) = (0,0);
		(Amult[30] => Cmult[15]) = (0,0);
		(Amult[31] => Cmult[15]) = (0,0);
		(Bmult[0]  => Cmult[15]) = (0,0);
		(Bmult[1]  => Cmult[15]) = (0,0);
		(Bmult[2]  => Cmult[15]) = (0,0);
		(Bmult[3]  => Cmult[15]) = (0,0);
		(Bmult[4]  => Cmult[15]) = (0,0);
		(Bmult[5]  => Cmult[15]) = (0,0);
		(Bmult[6]  => Cmult[15]) = (0,0);
		(Bmult[7]  => Cmult[15]) = (0,0);
		(Bmult[8]  => Cmult[15]) = (0,0);
		(Bmult[9]  => Cmult[15]) = (0,0);
		(Bmult[10] => Cmult[15]) = (0,0);
		(Bmult[11] => Cmult[15]) = (0,0);
		(Bmult[12] => Cmult[15]) = (0,0);
		(Bmult[13] => Cmult[15]) = (0,0);
		(Bmult[14] => Cmult[15]) = (0,0);
		(Bmult[15] => Cmult[15]) = (0,0);
		(Bmult[16] => Cmult[15]) = (0,0);
		(Bmult[17] => Cmult[15]) = (0,0);
		(Bmult[18] => Cmult[15]) = (0,0);
		(Bmult[19] => Cmult[15]) = (0,0);
		(Bmult[20] => Cmult[15]) = (0,0);
		(Bmult[21] => Cmult[15]) = (0,0);
		(Bmult[22] => Cmult[15]) = (0,0);
		(Bmult[23] => Cmult[15]) = (0,0);
		(Bmult[24] => Cmult[15]) = (0,0);
		(Bmult[25] => Cmult[15]) = (0,0);
		(Bmult[26] => Cmult[15]) = (0,0);
		(Bmult[27] => Cmult[15]) = (0,0);
		(Bmult[28] => Cmult[15]) = (0,0);
		(Bmult[29] => Cmult[15]) = (0,0);
		(Bmult[30] => Cmult[15]) = (0,0);
		(Bmult[31] => Cmult[15]) = (0,0);		
		(Valid_mult[0] => Cmult[15]) = (0,0);
		(Valid_mult[1] => Cmult[15]) = (0,0);
		(sel_mul_32x32 => Cmult[15]) = (0,0);
		(Amult[0]  => Cmult[16]) = (0,0);
		(Amult[1]  => Cmult[16]) = (0,0);
		(Amult[2]  => Cmult[16]) = (0,0);
		(Amult[3]  => Cmult[16]) = (0,0);
		(Amult[4]  => Cmult[16]) = (0,0);
		(Amult[5]  => Cmult[16]) = (0,0);
		(Amult[6]  => Cmult[16]) = (0,0);
		(Amult[7]  => Cmult[16]) = (0,0);
		(Amult[8]  => Cmult[16]) = (0,0);
		(Amult[9]  => Cmult[16]) = (0,0);
		(Amult[10] => Cmult[16]) = (0,0);
		(Amult[11] => Cmult[16]) = (0,0);
		(Amult[12] => Cmult[16]) = (0,0);
		(Amult[13] => Cmult[16]) = (0,0);
		(Amult[14] => Cmult[16]) = (0,0);
		(Amult[15] => Cmult[16]) = (0,0);
		(Amult[16] => Cmult[16]) = (0,0);
		(Amult[17] => Cmult[16]) = (0,0);
		(Amult[18] => Cmult[16]) = (0,0);
		(Amult[19] => Cmult[16]) = (0,0);
		(Amult[20] => Cmult[16]) = (0,0);
		(Amult[21] => Cmult[16]) = (0,0);
		(Amult[22] => Cmult[16]) = (0,0);
		(Amult[23] => Cmult[16]) = (0,0);
		(Amult[24] => Cmult[16]) = (0,0);
		(Amult[25] => Cmult[16]) = (0,0);
		(Amult[26] => Cmult[16]) = (0,0);
		(Amult[27] => Cmult[16]) = (0,0);
		(Amult[28] => Cmult[16]) = (0,0);
		(Amult[29] => Cmult[16]) = (0,0);
		(Amult[30] => Cmult[16]) = (0,0);
		(Amult[31] => Cmult[16]) = (0,0);
		(Bmult[0]  => Cmult[16]) = (0,0);
		(Bmult[1]  => Cmult[16]) = (0,0);
		(Bmult[2]  => Cmult[16]) = (0,0);
		(Bmult[3]  => Cmult[16]) = (0,0);
		(Bmult[4]  => Cmult[16]) = (0,0);
		(Bmult[5]  => Cmult[16]) = (0,0);
		(Bmult[6]  => Cmult[16]) = (0,0);
		(Bmult[7]  => Cmult[16]) = (0,0);
		(Bmult[8]  => Cmult[16]) = (0,0);
		(Bmult[9]  => Cmult[16]) = (0,0);
		(Bmult[10] => Cmult[16]) = (0,0);
		(Bmult[11] => Cmult[16]) = (0,0);
		(Bmult[12] => Cmult[16]) = (0,0);
		(Bmult[13] => Cmult[16]) = (0,0);
		(Bmult[14] => Cmult[16]) = (0,0);
		(Bmult[15] => Cmult[16]) = (0,0);
		(Bmult[16] => Cmult[16]) = (0,0);
		(Bmult[17] => Cmult[16]) = (0,0);
		(Bmult[18] => Cmult[16]) = (0,0);
		(Bmult[19] => Cmult[16]) = (0,0);
		(Bmult[20] => Cmult[16]) = (0,0);
		(Bmult[21] => Cmult[16]) = (0,0);
		(Bmult[22] => Cmult[16]) = (0,0);
		(Bmult[23] => Cmult[16]) = (0,0);
		(Bmult[24] => Cmult[16]) = (0,0);
		(Bmult[25] => Cmult[16]) = (0,0);
		(Bmult[26] => Cmult[16]) = (0,0);
		(Bmult[27] => Cmult[16]) = (0,0);
		(Bmult[28] => Cmult[16]) = (0,0);
		(Bmult[29] => Cmult[16]) = (0,0);
		(Bmult[30] => Cmult[16]) = (0,0);
		(Bmult[31] => Cmult[16]) = (0,0);		
		(Valid_mult[0] => Cmult[16]) = (0,0);
		(Valid_mult[1] => Cmult[16]) = (0,0);
		(sel_mul_32x32 => Cmult[16]) = (0,0);
		(Amult[0]  => Cmult[17]) = (0,0);
		(Amult[1]  => Cmult[17]) = (0,0);
		(Amult[2]  => Cmult[17]) = (0,0);
		(Amult[3]  => Cmult[17]) = (0,0);
		(Amult[4]  => Cmult[17]) = (0,0);
		(Amult[5]  => Cmult[17]) = (0,0);
		(Amult[6]  => Cmult[17]) = (0,0);
		(Amult[7]  => Cmult[17]) = (0,0);
		(Amult[8]  => Cmult[17]) = (0,0);
		(Amult[9]  => Cmult[17]) = (0,0);
		(Amult[10] => Cmult[17]) = (0,0);
		(Amult[11] => Cmult[17]) = (0,0);
		(Amult[12] => Cmult[17]) = (0,0);
		(Amult[13] => Cmult[17]) = (0,0);
		(Amult[14] => Cmult[17]) = (0,0);
		(Amult[15] => Cmult[17]) = (0,0);
		(Amult[16] => Cmult[17]) = (0,0);
		(Amult[17] => Cmult[17]) = (0,0);
		(Amult[18] => Cmult[17]) = (0,0);
		(Amult[19] => Cmult[17]) = (0,0);
		(Amult[20] => Cmult[17]) = (0,0);
		(Amult[21] => Cmult[17]) = (0,0);
		(Amult[22] => Cmult[17]) = (0,0);
		(Amult[23] => Cmult[17]) = (0,0);
		(Amult[24] => Cmult[17]) = (0,0);
		(Amult[25] => Cmult[17]) = (0,0);
		(Amult[26] => Cmult[17]) = (0,0);
		(Amult[27] => Cmult[17]) = (0,0);
		(Amult[28] => Cmult[17]) = (0,0);
		(Amult[29] => Cmult[17]) = (0,0);
		(Amult[30] => Cmult[17]) = (0,0);
		(Amult[31] => Cmult[17]) = (0,0);
		(Bmult[0]  => Cmult[17]) = (0,0);
		(Bmult[1]  => Cmult[17]) = (0,0);
		(Bmult[2]  => Cmult[17]) = (0,0);
		(Bmult[3]  => Cmult[17]) = (0,0);
		(Bmult[4]  => Cmult[17]) = (0,0);
		(Bmult[5]  => Cmult[17]) = (0,0);
		(Bmult[6]  => Cmult[17]) = (0,0);
		(Bmult[7]  => Cmult[17]) = (0,0);
		(Bmult[8]  => Cmult[17]) = (0,0);
		(Bmult[9]  => Cmult[17]) = (0,0);
		(Bmult[10] => Cmult[17]) = (0,0);
		(Bmult[11] => Cmult[17]) = (0,0);
		(Bmult[12] => Cmult[17]) = (0,0);
		(Bmult[13] => Cmult[17]) = (0,0);
		(Bmult[14] => Cmult[17]) = (0,0);
		(Bmult[15] => Cmult[17]) = (0,0);
		(Bmult[16] => Cmult[17]) = (0,0);
		(Bmult[17] => Cmult[17]) = (0,0);
		(Bmult[18] => Cmult[17]) = (0,0);
		(Bmult[19] => Cmult[17]) = (0,0);
		(Bmult[20] => Cmult[17]) = (0,0);
		(Bmult[21] => Cmult[17]) = (0,0);
		(Bmult[22] => Cmult[17]) = (0,0);
		(Bmult[23] => Cmult[17]) = (0,0);
		(Bmult[24] => Cmult[17]) = (0,0);
		(Bmult[25] => Cmult[17]) = (0,0);
		(Bmult[26] => Cmult[17]) = (0,0);
		(Bmult[27] => Cmult[17]) = (0,0);
		(Bmult[28] => Cmult[17]) = (0,0);
		(Bmult[29] => Cmult[17]) = (0,0);
		(Bmult[30] => Cmult[17]) = (0,0);
		(Bmult[31] => Cmult[17]) = (0,0);		
		(Valid_mult[0] => Cmult[17]) = (0,0);
		(Valid_mult[1] => Cmult[17]) = (0,0);
		(sel_mul_32x32 => Cmult[17]) = (0,0);
		(Amult[0]  => Cmult[18]) = (0,0);
		(Amult[1]  => Cmult[18]) = (0,0);
		(Amult[2]  => Cmult[18]) = (0,0);
		(Amult[3]  => Cmult[18]) = (0,0);
		(Amult[4]  => Cmult[18]) = (0,0);
		(Amult[5]  => Cmult[18]) = (0,0);
		(Amult[6]  => Cmult[18]) = (0,0);
		(Amult[7]  => Cmult[18]) = (0,0);
		(Amult[8]  => Cmult[18]) = (0,0);
		(Amult[9]  => Cmult[18]) = (0,0);
		(Amult[10] => Cmult[18]) = (0,0);
		(Amult[11] => Cmult[18]) = (0,0);
		(Amult[12] => Cmult[18]) = (0,0);
		(Amult[13] => Cmult[18]) = (0,0);
		(Amult[14] => Cmult[18]) = (0,0);
		(Amult[15] => Cmult[18]) = (0,0);
		(Amult[16] => Cmult[18]) = (0,0);
		(Amult[17] => Cmult[18]) = (0,0);
		(Amult[18] => Cmult[18]) = (0,0);
		(Amult[19] => Cmult[18]) = (0,0);
		(Amult[20] => Cmult[18]) = (0,0);
		(Amult[21] => Cmult[18]) = (0,0);
		(Amult[22] => Cmult[18]) = (0,0);
		(Amult[23] => Cmult[18]) = (0,0);
		(Amult[24] => Cmult[18]) = (0,0);
		(Amult[25] => Cmult[18]) = (0,0);
		(Amult[26] => Cmult[18]) = (0,0);
		(Amult[27] => Cmult[18]) = (0,0);
		(Amult[28] => Cmult[18]) = (0,0);
		(Amult[29] => Cmult[18]) = (0,0);
		(Amult[30] => Cmult[18]) = (0,0);
		(Amult[31] => Cmult[18]) = (0,0);
		(Bmult[0]  => Cmult[18]) = (0,0);
		(Bmult[1]  => Cmult[18]) = (0,0);
		(Bmult[2]  => Cmult[18]) = (0,0);
		(Bmult[3]  => Cmult[18]) = (0,0);
		(Bmult[4]  => Cmult[18]) = (0,0);
		(Bmult[5]  => Cmult[18]) = (0,0);
		(Bmult[6]  => Cmult[18]) = (0,0);
		(Bmult[7]  => Cmult[18]) = (0,0);
		(Bmult[8]  => Cmult[18]) = (0,0);
		(Bmult[9]  => Cmult[18]) = (0,0);
		(Bmult[10] => Cmult[18]) = (0,0);
		(Bmult[11] => Cmult[18]) = (0,0);
		(Bmult[12] => Cmult[18]) = (0,0);
		(Bmult[13] => Cmult[18]) = (0,0);
		(Bmult[14] => Cmult[18]) = (0,0);
		(Bmult[15] => Cmult[18]) = (0,0);
		(Bmult[16] => Cmult[18]) = (0,0);
		(Bmult[17] => Cmult[18]) = (0,0);
		(Bmult[18] => Cmult[18]) = (0,0);
		(Bmult[19] => Cmult[18]) = (0,0);
		(Bmult[20] => Cmult[18]) = (0,0);
		(Bmult[21] => Cmult[18]) = (0,0);
		(Bmult[22] => Cmult[18]) = (0,0);
		(Bmult[23] => Cmult[18]) = (0,0);
		(Bmult[24] => Cmult[18]) = (0,0);
		(Bmult[25] => Cmult[18]) = (0,0);
		(Bmult[26] => Cmult[18]) = (0,0);
		(Bmult[27] => Cmult[18]) = (0,0);
		(Bmult[28] => Cmult[18]) = (0,0);
		(Bmult[29] => Cmult[18]) = (0,0);
		(Bmult[30] => Cmult[18]) = (0,0);
		(Bmult[31] => Cmult[18]) = (0,0);		
		(Valid_mult[0] => Cmult[18]) = (0,0);
		(Valid_mult[1] => Cmult[18]) = (0,0);
		(sel_mul_32x32 => Cmult[18]) = (0,0);	
		(Amult[0]  => Cmult[19]) = (0,0);
		(Amult[1]  => Cmult[19]) = (0,0);
		(Amult[2]  => Cmult[19]) = (0,0);
		(Amult[3]  => Cmult[19]) = (0,0);
		(Amult[4]  => Cmult[19]) = (0,0);
		(Amult[5]  => Cmult[19]) = (0,0);
		(Amult[6]  => Cmult[19]) = (0,0);
		(Amult[7]  => Cmult[19]) = (0,0);
		(Amult[8]  => Cmult[19]) = (0,0);
		(Amult[9]  => Cmult[19]) = (0,0);
		(Amult[10] => Cmult[19]) = (0,0);
		(Amult[11] => Cmult[19]) = (0,0);
		(Amult[12] => Cmult[19]) = (0,0);
		(Amult[13] => Cmult[19]) = (0,0);
		(Amult[14] => Cmult[19]) = (0,0);
		(Amult[15] => Cmult[19]) = (0,0);
		(Amult[16] => Cmult[19]) = (0,0);
		(Amult[17] => Cmult[19]) = (0,0);
		(Amult[18] => Cmult[19]) = (0,0);
		(Amult[19] => Cmult[19]) = (0,0);
		(Amult[20] => Cmult[19]) = (0,0);
		(Amult[21] => Cmult[19]) = (0,0);
		(Amult[22] => Cmult[19]) = (0,0);
		(Amult[23] => Cmult[19]) = (0,0);
		(Amult[24] => Cmult[19]) = (0,0);
		(Amult[25] => Cmult[19]) = (0,0);
		(Amult[26] => Cmult[19]) = (0,0);
		(Amult[27] => Cmult[19]) = (0,0);
		(Amult[28] => Cmult[19]) = (0,0);
		(Amult[29] => Cmult[19]) = (0,0);
		(Amult[30] => Cmult[19]) = (0,0);
		(Amult[31] => Cmult[19]) = (0,0);
		(Bmult[0]  => Cmult[19]) = (0,0);
		(Bmult[1]  => Cmult[19]) = (0,0);
		(Bmult[2]  => Cmult[19]) = (0,0);
		(Bmult[3]  => Cmult[19]) = (0,0);
		(Bmult[4]  => Cmult[19]) = (0,0);
		(Bmult[5]  => Cmult[19]) = (0,0);
		(Bmult[6]  => Cmult[19]) = (0,0);
		(Bmult[7]  => Cmult[19]) = (0,0);
		(Bmult[8]  => Cmult[19]) = (0,0);
		(Bmult[9]  => Cmult[19]) = (0,0);
		(Bmult[10] => Cmult[19]) = (0,0);
		(Bmult[11] => Cmult[19]) = (0,0);
		(Bmult[12] => Cmult[19]) = (0,0);
		(Bmult[13] => Cmult[19]) = (0,0);
		(Bmult[14] => Cmult[19]) = (0,0);
		(Bmult[15] => Cmult[19]) = (0,0);
		(Bmult[16] => Cmult[19]) = (0,0);
		(Bmult[17] => Cmult[19]) = (0,0);
		(Bmult[18] => Cmult[19]) = (0,0);
		(Bmult[19] => Cmult[19]) = (0,0);
		(Bmult[20] => Cmult[19]) = (0,0);
		(Bmult[21] => Cmult[19]) = (0,0);
		(Bmult[22] => Cmult[19]) = (0,0);
		(Bmult[23] => Cmult[19]) = (0,0);
		(Bmult[24] => Cmult[19]) = (0,0);
		(Bmult[25] => Cmult[19]) = (0,0);
		(Bmult[26] => Cmult[19]) = (0,0);
		(Bmult[27] => Cmult[19]) = (0,0);
		(Bmult[28] => Cmult[19]) = (0,0);
		(Bmult[29] => Cmult[19]) = (0,0);
		(Bmult[30] => Cmult[19]) = (0,0);
		(Bmult[31] => Cmult[19]) = (0,0);		
		(Valid_mult[0] => Cmult[19]) = (0,0);
		(Valid_mult[1] => Cmult[19]) = (0,0);
		(sel_mul_32x32 => Cmult[19]) = (0,0);
		(Amult[0]  => Cmult[20]) = (0,0);
		(Amult[1]  => Cmult[20]) = (0,0);
		(Amult[2]  => Cmult[20]) = (0,0);
		(Amult[3]  => Cmult[20]) = (0,0);
		(Amult[4]  => Cmult[20]) = (0,0);
		(Amult[5]  => Cmult[20]) = (0,0);
		(Amult[6]  => Cmult[20]) = (0,0);
		(Amult[7]  => Cmult[20]) = (0,0);
		(Amult[8]  => Cmult[20]) = (0,0);
		(Amult[9]  => Cmult[20]) = (0,0);
		(Amult[10] => Cmult[20]) = (0,0);
		(Amult[11] => Cmult[20]) = (0,0);
		(Amult[12] => Cmult[20]) = (0,0);
		(Amult[13] => Cmult[20]) = (0,0);
		(Amult[14] => Cmult[20]) = (0,0);
		(Amult[15] => Cmult[20]) = (0,0);
		(Amult[16] => Cmult[20]) = (0,0);
		(Amult[17] => Cmult[20]) = (0,0);
		(Amult[18] => Cmult[20]) = (0,0);
		(Amult[19] => Cmult[20]) = (0,0);
		(Amult[20] => Cmult[20]) = (0,0);
		(Amult[21] => Cmult[20]) = (0,0);
		(Amult[22] => Cmult[20]) = (0,0);
		(Amult[23] => Cmult[20]) = (0,0);
		(Amult[24] => Cmult[20]) = (0,0);
		(Amult[25] => Cmult[20]) = (0,0);
		(Amult[26] => Cmult[20]) = (0,0);
		(Amult[27] => Cmult[20]) = (0,0);
		(Amult[28] => Cmult[20]) = (0,0);
		(Amult[29] => Cmult[20]) = (0,0);
		(Amult[30] => Cmult[20]) = (0,0);
		(Amult[31] => Cmult[20]) = (0,0);
		(Bmult[0]  => Cmult[20]) = (0,0);
		(Bmult[1]  => Cmult[20]) = (0,0);
		(Bmult[2]  => Cmult[20]) = (0,0);
		(Bmult[3]  => Cmult[20]) = (0,0);
		(Bmult[4]  => Cmult[20]) = (0,0);
		(Bmult[5]  => Cmult[20]) = (0,0);
		(Bmult[6]  => Cmult[20]) = (0,0);
		(Bmult[7]  => Cmult[20]) = (0,0);
		(Bmult[8]  => Cmult[20]) = (0,0);
		(Bmult[9]  => Cmult[20]) = (0,0);
		(Bmult[10] => Cmult[20]) = (0,0);
		(Bmult[11] => Cmult[20]) = (0,0);
		(Bmult[12] => Cmult[20]) = (0,0);
		(Bmult[13] => Cmult[20]) = (0,0);
		(Bmult[14] => Cmult[20]) = (0,0);
		(Bmult[15] => Cmult[20]) = (0,0);
		(Bmult[16] => Cmult[20]) = (0,0);
		(Bmult[17] => Cmult[20]) = (0,0);
		(Bmult[18] => Cmult[20]) = (0,0);
		(Bmult[19] => Cmult[20]) = (0,0);
		(Bmult[20] => Cmult[20]) = (0,0);
		(Bmult[21] => Cmult[20]) = (0,0);
		(Bmult[22] => Cmult[20]) = (0,0);
		(Bmult[23] => Cmult[20]) = (0,0);
		(Bmult[24] => Cmult[20]) = (0,0);
		(Bmult[25] => Cmult[20]) = (0,0);
		(Bmult[26] => Cmult[20]) = (0,0);
		(Bmult[27] => Cmult[20]) = (0,0);
		(Bmult[28] => Cmult[20]) = (0,0);
		(Bmult[29] => Cmult[20]) = (0,0);
		(Bmult[30] => Cmult[20]) = (0,0);
		(Bmult[31] => Cmult[20]) = (0,0);		
		(Valid_mult[0] => Cmult[20]) = (0,0);
		(Valid_mult[1] => Cmult[20]) = (0,0);
		(sel_mul_32x32 => Cmult[20]) = (0,0);
		(Amult[0]  => Cmult[21]) = (0,0);
		(Amult[1]  => Cmult[21]) = (0,0);
		(Amult[2]  => Cmult[21]) = (0,0);
		(Amult[3]  => Cmult[21]) = (0,0);
		(Amult[4]  => Cmult[21]) = (0,0);
		(Amult[5]  => Cmult[21]) = (0,0);
		(Amult[6]  => Cmult[21]) = (0,0);
		(Amult[7]  => Cmult[21]) = (0,0);
		(Amult[8]  => Cmult[21]) = (0,0);
		(Amult[9]  => Cmult[21]) = (0,0);
		(Amult[10] => Cmult[21]) = (0,0);
		(Amult[11] => Cmult[21]) = (0,0);
		(Amult[12] => Cmult[21]) = (0,0);
		(Amult[13] => Cmult[21]) = (0,0);
		(Amult[14] => Cmult[21]) = (0,0);
		(Amult[15] => Cmult[21]) = (0,0);
		(Amult[16] => Cmult[21]) = (0,0);
		(Amult[17] => Cmult[21]) = (0,0);
		(Amult[18] => Cmult[21]) = (0,0);
		(Amult[19] => Cmult[21]) = (0,0);
		(Amult[20] => Cmult[21]) = (0,0);
		(Amult[21] => Cmult[21]) = (0,0);
		(Amult[22] => Cmult[21]) = (0,0);
		(Amult[23] => Cmult[21]) = (0,0);
		(Amult[24] => Cmult[21]) = (0,0);
		(Amult[25] => Cmult[21]) = (0,0);
		(Amult[26] => Cmult[21]) = (0,0);
		(Amult[27] => Cmult[21]) = (0,0);
		(Amult[28] => Cmult[21]) = (0,0);
		(Amult[29] => Cmult[21]) = (0,0);
		(Amult[30] => Cmult[21]) = (0,0);
		(Amult[31] => Cmult[21]) = (0,0);
		(Bmult[0]  => Cmult[21]) = (0,0);
		(Bmult[1]  => Cmult[21]) = (0,0);
		(Bmult[2]  => Cmult[21]) = (0,0);
		(Bmult[3]  => Cmult[21]) = (0,0);
		(Bmult[4]  => Cmult[21]) = (0,0);
		(Bmult[5]  => Cmult[21]) = (0,0);
		(Bmult[6]  => Cmult[21]) = (0,0);
		(Bmult[7]  => Cmult[21]) = (0,0);
		(Bmult[8]  => Cmult[21]) = (0,0);
		(Bmult[9]  => Cmult[21]) = (0,0);
		(Bmult[10] => Cmult[21]) = (0,0);
		(Bmult[11] => Cmult[21]) = (0,0);
		(Bmult[12] => Cmult[21]) = (0,0);
		(Bmult[13] => Cmult[21]) = (0,0);
		(Bmult[14] => Cmult[21]) = (0,0);
		(Bmult[15] => Cmult[21]) = (0,0);
		(Bmult[16] => Cmult[21]) = (0,0);
		(Bmult[17] => Cmult[21]) = (0,0);
		(Bmult[18] => Cmult[21]) = (0,0);
		(Bmult[19] => Cmult[21]) = (0,0);
		(Bmult[20] => Cmult[21]) = (0,0);
		(Bmult[21] => Cmult[21]) = (0,0);
		(Bmult[22] => Cmult[21]) = (0,0);
		(Bmult[23] => Cmult[21]) = (0,0);
		(Bmult[24] => Cmult[21]) = (0,0);
		(Bmult[25] => Cmult[21]) = (0,0);
		(Bmult[26] => Cmult[21]) = (0,0);
		(Bmult[27] => Cmult[21]) = (0,0);
		(Bmult[28] => Cmult[21]) = (0,0);
		(Bmult[29] => Cmult[21]) = (0,0);
		(Bmult[30] => Cmult[21]) = (0,0);
		(Bmult[31] => Cmult[21]) = (0,0);		
		(Valid_mult[0] => Cmult[21]) = (0,0);
		(Valid_mult[1] => Cmult[21]) = (0,0);
		(sel_mul_32x32 => Cmult[21]) = (0,0);
		(Amult[0]  => Cmult[22]) = (0,0);
		(Amult[1]  => Cmult[22]) = (0,0);
		(Amult[2]  => Cmult[22]) = (0,0);
		(Amult[3]  => Cmult[22]) = (0,0);
		(Amult[4]  => Cmult[22]) = (0,0);
		(Amult[5]  => Cmult[22]) = (0,0);
		(Amult[6]  => Cmult[22]) = (0,0);
		(Amult[7]  => Cmult[22]) = (0,0);
		(Amult[8]  => Cmult[22]) = (0,0);
		(Amult[9]  => Cmult[22]) = (0,0);
		(Amult[10] => Cmult[22]) = (0,0);
		(Amult[11] => Cmult[22]) = (0,0);
		(Amult[12] => Cmult[22]) = (0,0);
		(Amult[13] => Cmult[22]) = (0,0);
		(Amult[14] => Cmult[22]) = (0,0);
		(Amult[15] => Cmult[22]) = (0,0);
		(Amult[16] => Cmult[22]) = (0,0);
		(Amult[17] => Cmult[22]) = (0,0);
		(Amult[18] => Cmult[22]) = (0,0);
		(Amult[19] => Cmult[22]) = (0,0);
		(Amult[20] => Cmult[22]) = (0,0);
		(Amult[21] => Cmult[22]) = (0,0);
		(Amult[22] => Cmult[22]) = (0,0);
		(Amult[23] => Cmult[22]) = (0,0);
		(Amult[24] => Cmult[22]) = (0,0);
		(Amult[25] => Cmult[22]) = (0,0);
		(Amult[26] => Cmult[22]) = (0,0);
		(Amult[27] => Cmult[22]) = (0,0);
		(Amult[28] => Cmult[22]) = (0,0);
		(Amult[29] => Cmult[22]) = (0,0);
		(Amult[30] => Cmult[22]) = (0,0);
		(Amult[31] => Cmult[22]) = (0,0);
		(Bmult[0]  => Cmult[22]) = (0,0);
		(Bmult[1]  => Cmult[22]) = (0,0);
		(Bmult[2]  => Cmult[22]) = (0,0);
		(Bmult[3]  => Cmult[22]) = (0,0);
		(Bmult[4]  => Cmult[22]) = (0,0);
		(Bmult[5]  => Cmult[22]) = (0,0);
		(Bmult[6]  => Cmult[22]) = (0,0);
		(Bmult[7]  => Cmult[22]) = (0,0);
		(Bmult[8]  => Cmult[22]) = (0,0);
		(Bmult[9]  => Cmult[22]) = (0,0);
		(Bmult[10] => Cmult[22]) = (0,0);
		(Bmult[11] => Cmult[22]) = (0,0);
		(Bmult[12] => Cmult[22]) = (0,0);
		(Bmult[13] => Cmult[22]) = (0,0);
		(Bmult[14] => Cmult[22]) = (0,0);
		(Bmult[15] => Cmult[22]) = (0,0);
		(Bmult[16] => Cmult[22]) = (0,0);
		(Bmult[17] => Cmult[22]) = (0,0);
		(Bmult[18] => Cmult[22]) = (0,0);
		(Bmult[19] => Cmult[22]) = (0,0);
		(Bmult[20] => Cmult[22]) = (0,0);
		(Bmult[21] => Cmult[22]) = (0,0);
		(Bmult[22] => Cmult[22]) = (0,0);
		(Bmult[23] => Cmult[22]) = (0,0);
		(Bmult[24] => Cmult[22]) = (0,0);
		(Bmult[25] => Cmult[22]) = (0,0);
		(Bmult[26] => Cmult[22]) = (0,0);
		(Bmult[27] => Cmult[22]) = (0,0);
		(Bmult[28] => Cmult[22]) = (0,0);
		(Bmult[29] => Cmult[22]) = (0,0);
		(Bmult[30] => Cmult[22]) = (0,0);
		(Bmult[31] => Cmult[22]) = (0,0);		
		(Valid_mult[0] => Cmult[22]) = (0,0);
		(Valid_mult[1] => Cmult[22]) = (0,0);
		(sel_mul_32x32 => Cmult[22]) = (0,0);
		(Amult[0]  => Cmult[23]) = (0,0);
		(Amult[1]  => Cmult[23]) = (0,0);
		(Amult[2]  => Cmult[23]) = (0,0);
		(Amult[3]  => Cmult[23]) = (0,0);
		(Amult[4]  => Cmult[23]) = (0,0);
		(Amult[5]  => Cmult[23]) = (0,0);
		(Amult[6]  => Cmult[23]) = (0,0);
		(Amult[7]  => Cmult[23]) = (0,0);
		(Amult[8]  => Cmult[23]) = (0,0);
		(Amult[9]  => Cmult[23]) = (0,0);
		(Amult[10] => Cmult[23]) = (0,0);
		(Amult[11] => Cmult[23]) = (0,0);
		(Amult[12] => Cmult[23]) = (0,0);
		(Amult[13] => Cmult[23]) = (0,0);
		(Amult[14] => Cmult[23]) = (0,0);
		(Amult[15] => Cmult[23]) = (0,0);
		(Amult[16] => Cmult[23]) = (0,0);
		(Amult[17] => Cmult[23]) = (0,0);
		(Amult[18] => Cmult[23]) = (0,0);
		(Amult[19] => Cmult[23]) = (0,0);
		(Amult[20] => Cmult[23]) = (0,0);
		(Amult[21] => Cmult[23]) = (0,0);
		(Amult[22] => Cmult[23]) = (0,0);
		(Amult[23] => Cmult[23]) = (0,0);
		(Amult[24] => Cmult[23]) = (0,0);
		(Amult[25] => Cmult[23]) = (0,0);
		(Amult[26] => Cmult[23]) = (0,0);
		(Amult[27] => Cmult[23]) = (0,0);
		(Amult[28] => Cmult[23]) = (0,0);
		(Amult[29] => Cmult[23]) = (0,0);
		(Amult[30] => Cmult[23]) = (0,0);
		(Amult[31] => Cmult[23]) = (0,0);
		(Bmult[0]  => Cmult[23]) = (0,0);
		(Bmult[1]  => Cmult[23]) = (0,0);
		(Bmult[2]  => Cmult[23]) = (0,0);
		(Bmult[3]  => Cmult[23]) = (0,0);
		(Bmult[4]  => Cmult[23]) = (0,0);
		(Bmult[5]  => Cmult[23]) = (0,0);
		(Bmult[6]  => Cmult[23]) = (0,0);
		(Bmult[7]  => Cmult[23]) = (0,0);
		(Bmult[8]  => Cmult[23]) = (0,0);
		(Bmult[9]  => Cmult[23]) = (0,0);
		(Bmult[10] => Cmult[23]) = (0,0);
		(Bmult[11] => Cmult[23]) = (0,0);
		(Bmult[12] => Cmult[23]) = (0,0);
		(Bmult[13] => Cmult[23]) = (0,0);
		(Bmult[14] => Cmult[23]) = (0,0);
		(Bmult[15] => Cmult[23]) = (0,0);
		(Bmult[16] => Cmult[23]) = (0,0);
		(Bmult[17] => Cmult[23]) = (0,0);
		(Bmult[18] => Cmult[23]) = (0,0);
		(Bmult[19] => Cmult[23]) = (0,0);
		(Bmult[20] => Cmult[23]) = (0,0);
		(Bmult[21] => Cmult[23]) = (0,0);
		(Bmult[22] => Cmult[23]) = (0,0);
		(Bmult[23] => Cmult[23]) = (0,0);
		(Bmult[24] => Cmult[23]) = (0,0);
		(Bmult[25] => Cmult[23]) = (0,0);
		(Bmult[26] => Cmult[23]) = (0,0);
		(Bmult[27] => Cmult[23]) = (0,0);
		(Bmult[28] => Cmult[23]) = (0,0);
		(Bmult[29] => Cmult[23]) = (0,0);
		(Bmult[30] => Cmult[23]) = (0,0);
		(Bmult[31] => Cmult[23]) = (0,0);		
		(Valid_mult[0] => Cmult[23]) = (0,0);
		(Valid_mult[1] => Cmult[23]) = (0,0);
		(sel_mul_32x32 => Cmult[23]) = (0,0);
		(Amult[0]  => Cmult[24]) = (0,0);
		(Amult[1]  => Cmult[24]) = (0,0);
		(Amult[2]  => Cmult[24]) = (0,0);
		(Amult[3]  => Cmult[24]) = (0,0);
		(Amult[4]  => Cmult[24]) = (0,0);
		(Amult[5]  => Cmult[24]) = (0,0);
		(Amult[6]  => Cmult[24]) = (0,0);
		(Amult[7]  => Cmult[24]) = (0,0);
		(Amult[8]  => Cmult[24]) = (0,0);
		(Amult[9]  => Cmult[24]) = (0,0);
		(Amult[10] => Cmult[24]) = (0,0);
		(Amult[11] => Cmult[24]) = (0,0);
		(Amult[12] => Cmult[24]) = (0,0);
		(Amult[13] => Cmult[24]) = (0,0);
		(Amult[14] => Cmult[24]) = (0,0);
		(Amult[15] => Cmult[24]) = (0,0);
		(Amult[16] => Cmult[24]) = (0,0);
		(Amult[17] => Cmult[24]) = (0,0);
		(Amult[18] => Cmult[24]) = (0,0);
		(Amult[19] => Cmult[24]) = (0,0);
		(Amult[20] => Cmult[24]) = (0,0);
		(Amult[21] => Cmult[24]) = (0,0);
		(Amult[22] => Cmult[24]) = (0,0);
		(Amult[23] => Cmult[24]) = (0,0);
		(Amult[24] => Cmult[24]) = (0,0);
		(Amult[25] => Cmult[24]) = (0,0);
		(Amult[26] => Cmult[24]) = (0,0);
		(Amult[27] => Cmult[24]) = (0,0);
		(Amult[28] => Cmult[24]) = (0,0);
		(Amult[29] => Cmult[24]) = (0,0);
		(Amult[30] => Cmult[24]) = (0,0);
		(Amult[31] => Cmult[24]) = (0,0);
		(Bmult[0]  => Cmult[24]) = (0,0);
		(Bmult[1]  => Cmult[24]) = (0,0);
		(Bmult[2]  => Cmult[24]) = (0,0);
		(Bmult[3]  => Cmult[24]) = (0,0);
		(Bmult[4]  => Cmult[24]) = (0,0);
		(Bmult[5]  => Cmult[24]) = (0,0);
		(Bmult[6]  => Cmult[24]) = (0,0);
		(Bmult[7]  => Cmult[24]) = (0,0);
		(Bmult[8]  => Cmult[24]) = (0,0);
		(Bmult[9]  => Cmult[24]) = (0,0);
		(Bmult[10] => Cmult[24]) = (0,0);
		(Bmult[11] => Cmult[24]) = (0,0);
		(Bmult[12] => Cmult[24]) = (0,0);
		(Bmult[13] => Cmult[24]) = (0,0);
		(Bmult[14] => Cmult[24]) = (0,0);
		(Bmult[15] => Cmult[24]) = (0,0);
		(Bmult[16] => Cmult[24]) = (0,0);
		(Bmult[17] => Cmult[24]) = (0,0);
		(Bmult[18] => Cmult[24]) = (0,0);
		(Bmult[19] => Cmult[24]) = (0,0);
		(Bmult[20] => Cmult[24]) = (0,0);
		(Bmult[21] => Cmult[24]) = (0,0);
		(Bmult[22] => Cmult[24]) = (0,0);
		(Bmult[23] => Cmult[24]) = (0,0);
		(Bmult[24] => Cmult[24]) = (0,0);
		(Bmult[25] => Cmult[24]) = (0,0);
		(Bmult[26] => Cmult[24]) = (0,0);
		(Bmult[27] => Cmult[24]) = (0,0);
		(Bmult[28] => Cmult[24]) = (0,0);
		(Bmult[29] => Cmult[24]) = (0,0);
		(Bmult[30] => Cmult[24]) = (0,0);
		(Bmult[31] => Cmult[24]) = (0,0);		
		(Valid_mult[0] => Cmult[24]) = (0,0);
		(Valid_mult[1] => Cmult[24]) = (0,0);
		(sel_mul_32x32 => Cmult[24]) = (0,0);
		(Amult[0]  => Cmult[25]) = (0,0);
		(Amult[1]  => Cmult[25]) = (0,0);
		(Amult[2]  => Cmult[25]) = (0,0);
		(Amult[3]  => Cmult[25]) = (0,0);
		(Amult[4]  => Cmult[25]) = (0,0);
		(Amult[5]  => Cmult[25]) = (0,0);
		(Amult[6]  => Cmult[25]) = (0,0);
		(Amult[7]  => Cmult[25]) = (0,0);
		(Amult[8]  => Cmult[25]) = (0,0);
		(Amult[9]  => Cmult[25]) = (0,0);
		(Amult[10] => Cmult[25]) = (0,0);
		(Amult[11] => Cmult[25]) = (0,0);
		(Amult[12] => Cmult[25]) = (0,0);
		(Amult[13] => Cmult[25]) = (0,0);
		(Amult[14] => Cmult[25]) = (0,0);
		(Amult[15] => Cmult[25]) = (0,0);
		(Amult[16] => Cmult[25]) = (0,0);
		(Amult[17] => Cmult[25]) = (0,0);
		(Amult[18] => Cmult[25]) = (0,0);
		(Amult[19] => Cmult[25]) = (0,0);
		(Amult[20] => Cmult[25]) = (0,0);
		(Amult[21] => Cmult[25]) = (0,0);
		(Amult[22] => Cmult[25]) = (0,0);
		(Amult[23] => Cmult[25]) = (0,0);
		(Amult[24] => Cmult[25]) = (0,0);
		(Amult[25] => Cmult[25]) = (0,0);
		(Amult[26] => Cmult[25]) = (0,0);
		(Amult[27] => Cmult[25]) = (0,0);
		(Amult[28] => Cmult[25]) = (0,0);
		(Amult[29] => Cmult[25]) = (0,0);
		(Amult[30] => Cmult[25]) = (0,0);
		(Amult[31] => Cmult[25]) = (0,0);
		(Bmult[0]  => Cmult[25]) = (0,0);
		(Bmult[1]  => Cmult[25]) = (0,0);
		(Bmult[2]  => Cmult[25]) = (0,0);
		(Bmult[3]  => Cmult[25]) = (0,0);
		(Bmult[4]  => Cmult[25]) = (0,0);
		(Bmult[5]  => Cmult[25]) = (0,0);
		(Bmult[6]  => Cmult[25]) = (0,0);
		(Bmult[7]  => Cmult[25]) = (0,0);
		(Bmult[8]  => Cmult[25]) = (0,0);
		(Bmult[9]  => Cmult[25]) = (0,0);
		(Bmult[10] => Cmult[25]) = (0,0);
		(Bmult[11] => Cmult[25]) = (0,0);
		(Bmult[12] => Cmult[25]) = (0,0);
		(Bmult[13] => Cmult[25]) = (0,0);
		(Bmult[14] => Cmult[25]) = (0,0);
		(Bmult[15] => Cmult[25]) = (0,0);
		(Bmult[16] => Cmult[25]) = (0,0);
		(Bmult[17] => Cmult[25]) = (0,0);
		(Bmult[18] => Cmult[25]) = (0,0);
		(Bmult[19] => Cmult[25]) = (0,0);
		(Bmult[20] => Cmult[25]) = (0,0);
		(Bmult[21] => Cmult[25]) = (0,0);
		(Bmult[22] => Cmult[25]) = (0,0);
		(Bmult[23] => Cmult[25]) = (0,0);
		(Bmult[24] => Cmult[25]) = (0,0);
		(Bmult[25] => Cmult[25]) = (0,0);
		(Bmult[26] => Cmult[25]) = (0,0);
		(Bmult[27] => Cmult[25]) = (0,0);
		(Bmult[28] => Cmult[25]) = (0,0);
		(Bmult[29] => Cmult[25]) = (0,0);
		(Bmult[30] => Cmult[25]) = (0,0);
		(Bmult[31] => Cmult[25]) = (0,0);		
		(Valid_mult[0] => Cmult[25]) = (0,0);
		(Valid_mult[1] => Cmult[25]) = (0,0);
		(sel_mul_32x32 => Cmult[25]) = (0,0);
		(Amult[0]  => Cmult[26]) = (0,0);
		(Amult[1]  => Cmult[26]) = (0,0);
		(Amult[2]  => Cmult[26]) = (0,0);
		(Amult[3]  => Cmult[26]) = (0,0);
		(Amult[4]  => Cmult[26]) = (0,0);
		(Amult[5]  => Cmult[26]) = (0,0);
		(Amult[6]  => Cmult[26]) = (0,0);
		(Amult[7]  => Cmult[26]) = (0,0);
		(Amult[8]  => Cmult[26]) = (0,0);
		(Amult[9]  => Cmult[26]) = (0,0);
		(Amult[10] => Cmult[26]) = (0,0);
		(Amult[11] => Cmult[26]) = (0,0);
		(Amult[12] => Cmult[26]) = (0,0);
		(Amult[13] => Cmult[26]) = (0,0);
		(Amult[14] => Cmult[26]) = (0,0);
		(Amult[15] => Cmult[26]) = (0,0);
		(Amult[16] => Cmult[26]) = (0,0);
		(Amult[17] => Cmult[26]) = (0,0);
		(Amult[18] => Cmult[26]) = (0,0);
		(Amult[19] => Cmult[26]) = (0,0);
		(Amult[20] => Cmult[26]) = (0,0);
		(Amult[21] => Cmult[26]) = (0,0);
		(Amult[22] => Cmult[26]) = (0,0);
		(Amult[23] => Cmult[26]) = (0,0);
		(Amult[24] => Cmult[26]) = (0,0);
		(Amult[25] => Cmult[26]) = (0,0);
		(Amult[26] => Cmult[26]) = (0,0);
		(Amult[27] => Cmult[26]) = (0,0);
		(Amult[28] => Cmult[26]) = (0,0);
		(Amult[29] => Cmult[26]) = (0,0);
		(Amult[30] => Cmult[26]) = (0,0);
		(Amult[31] => Cmult[26]) = (0,0);
		(Bmult[0]  => Cmult[26]) = (0,0);
		(Bmult[1]  => Cmult[26]) = (0,0);
		(Bmult[2]  => Cmult[26]) = (0,0);
		(Bmult[3]  => Cmult[26]) = (0,0);
		(Bmult[4]  => Cmult[26]) = (0,0);
		(Bmult[5]  => Cmult[26]) = (0,0);
		(Bmult[6]  => Cmult[26]) = (0,0);
		(Bmult[7]  => Cmult[26]) = (0,0);
		(Bmult[8]  => Cmult[26]) = (0,0);
		(Bmult[9]  => Cmult[26]) = (0,0);
		(Bmult[10] => Cmult[26]) = (0,0);
		(Bmult[11] => Cmult[26]) = (0,0);
		(Bmult[12] => Cmult[26]) = (0,0);
		(Bmult[13] => Cmult[26]) = (0,0);
		(Bmult[14] => Cmult[26]) = (0,0);
		(Bmult[15] => Cmult[26]) = (0,0);
		(Bmult[16] => Cmult[26]) = (0,0);
		(Bmult[17] => Cmult[26]) = (0,0);
		(Bmult[18] => Cmult[26]) = (0,0);
		(Bmult[19] => Cmult[26]) = (0,0);
		(Bmult[20] => Cmult[26]) = (0,0);
		(Bmult[21] => Cmult[26]) = (0,0);
		(Bmult[22] => Cmult[26]) = (0,0);
		(Bmult[23] => Cmult[26]) = (0,0);
		(Bmult[24] => Cmult[26]) = (0,0);
		(Bmult[25] => Cmult[26]) = (0,0);
		(Bmult[26] => Cmult[26]) = (0,0);
		(Bmult[27] => Cmult[26]) = (0,0);
		(Bmult[28] => Cmult[26]) = (0,0);
		(Bmult[29] => Cmult[26]) = (0,0);
		(Bmult[30] => Cmult[26]) = (0,0);
		(Bmult[31] => Cmult[26]) = (0,0);		
		(Valid_mult[0] => Cmult[26]) = (0,0);
		(Valid_mult[1] => Cmult[26]) = (0,0);
		(sel_mul_32x32 => Cmult[26]) = (0,0);
		(Amult[0]  => Cmult[27]) = (0,0);
		(Amult[1]  => Cmult[27]) = (0,0);
		(Amult[2]  => Cmult[27]) = (0,0);
		(Amult[3]  => Cmult[27]) = (0,0);
		(Amult[4]  => Cmult[27]) = (0,0);
		(Amult[5]  => Cmult[27]) = (0,0);
		(Amult[6]  => Cmult[27]) = (0,0);
		(Amult[7]  => Cmult[27]) = (0,0);
		(Amult[8]  => Cmult[27]) = (0,0);
		(Amult[9]  => Cmult[27]) = (0,0);
		(Amult[10] => Cmult[27]) = (0,0);
		(Amult[11] => Cmult[27]) = (0,0);
		(Amult[12] => Cmult[27]) = (0,0);
		(Amult[13] => Cmult[27]) = (0,0);
		(Amult[14] => Cmult[27]) = (0,0);
		(Amult[15] => Cmult[27]) = (0,0);
		(Amult[16] => Cmult[27]) = (0,0);
		(Amult[17] => Cmult[27]) = (0,0);
		(Amult[18] => Cmult[27]) = (0,0);
		(Amult[19] => Cmult[27]) = (0,0);
		(Amult[20] => Cmult[27]) = (0,0);
		(Amult[21] => Cmult[27]) = (0,0);
		(Amult[22] => Cmult[27]) = (0,0);
		(Amult[23] => Cmult[27]) = (0,0);
		(Amult[24] => Cmult[27]) = (0,0);
		(Amult[25] => Cmult[27]) = (0,0);
		(Amult[26] => Cmult[27]) = (0,0);
		(Amult[27] => Cmult[27]) = (0,0);
		(Amult[28] => Cmult[27]) = (0,0);
		(Amult[29] => Cmult[27]) = (0,0);
		(Amult[30] => Cmult[27]) = (0,0);
		(Amult[31] => Cmult[27]) = (0,0);
		(Bmult[0]  => Cmult[27]) = (0,0);
		(Bmult[1]  => Cmult[27]) = (0,0);
		(Bmult[2]  => Cmult[27]) = (0,0);
		(Bmult[3]  => Cmult[27]) = (0,0);
		(Bmult[4]  => Cmult[27]) = (0,0);
		(Bmult[5]  => Cmult[27]) = (0,0);
		(Bmult[6]  => Cmult[27]) = (0,0);
		(Bmult[7]  => Cmult[27]) = (0,0);
		(Bmult[8]  => Cmult[27]) = (0,0);
		(Bmult[9]  => Cmult[27]) = (0,0);
		(Bmult[10] => Cmult[27]) = (0,0);
		(Bmult[11] => Cmult[27]) = (0,0);
		(Bmult[12] => Cmult[27]) = (0,0);
		(Bmult[13] => Cmult[27]) = (0,0);
		(Bmult[14] => Cmult[27]) = (0,0);
		(Bmult[15] => Cmult[27]) = (0,0);
		(Bmult[16] => Cmult[27]) = (0,0);
		(Bmult[17] => Cmult[27]) = (0,0);
		(Bmult[18] => Cmult[27]) = (0,0);
		(Bmult[19] => Cmult[27]) = (0,0);
		(Bmult[20] => Cmult[27]) = (0,0);
		(Bmult[21] => Cmult[27]) = (0,0);
		(Bmult[22] => Cmult[27]) = (0,0);
		(Bmult[23] => Cmult[27]) = (0,0);
		(Bmult[24] => Cmult[27]) = (0,0);
		(Bmult[25] => Cmult[27]) = (0,0);
		(Bmult[26] => Cmult[27]) = (0,0);
		(Bmult[27] => Cmult[27]) = (0,0);
		(Bmult[28] => Cmult[27]) = (0,0);
		(Bmult[29] => Cmult[27]) = (0,0);
		(Bmult[30] => Cmult[27]) = (0,0);
		(Bmult[31] => Cmult[27]) = (0,0);		
		(Valid_mult[0] => Cmult[27]) = (0,0);
		(Valid_mult[1] => Cmult[27]) = (0,0);
		(sel_mul_32x32 => Cmult[27]) = (0,0);
		(Amult[0]  => Cmult[28]) = (0,0);
		(Amult[1]  => Cmult[28]) = (0,0);
		(Amult[2]  => Cmult[28]) = (0,0);
		(Amult[3]  => Cmult[28]) = (0,0);
		(Amult[4]  => Cmult[28]) = (0,0);
		(Amult[5]  => Cmult[28]) = (0,0);
		(Amult[6]  => Cmult[28]) = (0,0);
		(Amult[7]  => Cmult[28]) = (0,0);
		(Amult[8]  => Cmult[28]) = (0,0);
		(Amult[9]  => Cmult[28]) = (0,0);
		(Amult[10] => Cmult[28]) = (0,0);
		(Amult[11] => Cmult[28]) = (0,0);
		(Amult[12] => Cmult[28]) = (0,0);
		(Amult[13] => Cmult[28]) = (0,0);
		(Amult[14] => Cmult[28]) = (0,0);
		(Amult[15] => Cmult[28]) = (0,0);
		(Amult[16] => Cmult[28]) = (0,0);
		(Amult[17] => Cmult[28]) = (0,0);
		(Amult[18] => Cmult[28]) = (0,0);
		(Amult[19] => Cmult[28]) = (0,0);
		(Amult[20] => Cmult[28]) = (0,0);
		(Amult[21] => Cmult[28]) = (0,0);
		(Amult[22] => Cmult[28]) = (0,0);
		(Amult[23] => Cmult[28]) = (0,0);
		(Amult[24] => Cmult[28]) = (0,0);
		(Amult[25] => Cmult[28]) = (0,0);
		(Amult[26] => Cmult[28]) = (0,0);
		(Amult[27] => Cmult[28]) = (0,0);
		(Amult[28] => Cmult[28]) = (0,0);
		(Amult[29] => Cmult[28]) = (0,0);
		(Amult[30] => Cmult[28]) = (0,0);
		(Amult[31] => Cmult[28]) = (0,0);
		(Bmult[0]  => Cmult[28]) = (0,0);
		(Bmult[1]  => Cmult[28]) = (0,0);
		(Bmult[2]  => Cmult[28]) = (0,0);
		(Bmult[3]  => Cmult[28]) = (0,0);
		(Bmult[4]  => Cmult[28]) = (0,0);
		(Bmult[5]  => Cmult[28]) = (0,0);
		(Bmult[6]  => Cmult[28]) = (0,0);
		(Bmult[7]  => Cmult[28]) = (0,0);
		(Bmult[8]  => Cmult[28]) = (0,0);
		(Bmult[9]  => Cmult[28]) = (0,0);
		(Bmult[10] => Cmult[28]) = (0,0);
		(Bmult[11] => Cmult[28]) = (0,0);
		(Bmult[12] => Cmult[28]) = (0,0);
		(Bmult[13] => Cmult[28]) = (0,0);
		(Bmult[14] => Cmult[28]) = (0,0);
		(Bmult[15] => Cmult[28]) = (0,0);
		(Bmult[16] => Cmult[28]) = (0,0);
		(Bmult[17] => Cmult[28]) = (0,0);
		(Bmult[18] => Cmult[28]) = (0,0);
		(Bmult[19] => Cmult[28]) = (0,0);
		(Bmult[20] => Cmult[28]) = (0,0);
		(Bmult[21] => Cmult[28]) = (0,0);
		(Bmult[22] => Cmult[28]) = (0,0);
		(Bmult[23] => Cmult[28]) = (0,0);
		(Bmult[24] => Cmult[28]) = (0,0);
		(Bmult[25] => Cmult[28]) = (0,0);
		(Bmult[26] => Cmult[28]) = (0,0);
		(Bmult[27] => Cmult[28]) = (0,0);
		(Bmult[28] => Cmult[28]) = (0,0);
		(Bmult[29] => Cmult[28]) = (0,0);
		(Bmult[30] => Cmult[28]) = (0,0);
		(Bmult[31] => Cmult[28]) = (0,0);		
		(Valid_mult[0] => Cmult[28]) = (0,0);
		(Valid_mult[1] => Cmult[28]) = (0,0);
		(sel_mul_32x32 => Cmult[28]) = (0,0);	
		(Amult[0]  => Cmult[29]) = (0,0);
		(Amult[1]  => Cmult[29]) = (0,0);
		(Amult[2]  => Cmult[29]) = (0,0);
		(Amult[3]  => Cmult[29]) = (0,0);
		(Amult[4]  => Cmult[29]) = (0,0);
		(Amult[5]  => Cmult[29]) = (0,0);
		(Amult[6]  => Cmult[29]) = (0,0);
		(Amult[7]  => Cmult[29]) = (0,0);
		(Amult[8]  => Cmult[29]) = (0,0);
		(Amult[9]  => Cmult[29]) = (0,0);
		(Amult[10] => Cmult[29]) = (0,0);
		(Amult[11] => Cmult[29]) = (0,0);
		(Amult[12] => Cmult[29]) = (0,0);
		(Amult[13] => Cmult[29]) = (0,0);
		(Amult[14] => Cmult[29]) = (0,0);
		(Amult[15] => Cmult[29]) = (0,0);
		(Amult[16] => Cmult[29]) = (0,0);
		(Amult[17] => Cmult[29]) = (0,0);
		(Amult[18] => Cmult[29]) = (0,0);
		(Amult[19] => Cmult[29]) = (0,0);
		(Amult[20] => Cmult[29]) = (0,0);
		(Amult[21] => Cmult[29]) = (0,0);
		(Amult[22] => Cmult[29]) = (0,0);
		(Amult[23] => Cmult[29]) = (0,0);
		(Amult[24] => Cmult[29]) = (0,0);
		(Amult[25] => Cmult[29]) = (0,0);
		(Amult[26] => Cmult[29]) = (0,0);
		(Amult[27] => Cmult[29]) = (0,0);
		(Amult[28] => Cmult[29]) = (0,0);
		(Amult[29] => Cmult[29]) = (0,0);
		(Amult[30] => Cmult[29]) = (0,0);
		(Amult[31] => Cmult[29]) = (0,0);
		(Bmult[0]  => Cmult[29]) = (0,0);
		(Bmult[1]  => Cmult[29]) = (0,0);
		(Bmult[2]  => Cmult[29]) = (0,0);
		(Bmult[3]  => Cmult[29]) = (0,0);
		(Bmult[4]  => Cmult[29]) = (0,0);
		(Bmult[5]  => Cmult[29]) = (0,0);
		(Bmult[6]  => Cmult[29]) = (0,0);
		(Bmult[7]  => Cmult[29]) = (0,0);
		(Bmult[8]  => Cmult[29]) = (0,0);
		(Bmult[9]  => Cmult[29]) = (0,0);
		(Bmult[10] => Cmult[29]) = (0,0);
		(Bmult[11] => Cmult[29]) = (0,0);
		(Bmult[12] => Cmult[29]) = (0,0);
		(Bmult[13] => Cmult[29]) = (0,0);
		(Bmult[14] => Cmult[29]) = (0,0);
		(Bmult[15] => Cmult[29]) = (0,0);
		(Bmult[16] => Cmult[29]) = (0,0);
		(Bmult[17] => Cmult[29]) = (0,0);
		(Bmult[18] => Cmult[29]) = (0,0);
		(Bmult[19] => Cmult[29]) = (0,0);
		(Bmult[20] => Cmult[29]) = (0,0);
		(Bmult[21] => Cmult[29]) = (0,0);
		(Bmult[22] => Cmult[29]) = (0,0);
		(Bmult[23] => Cmult[29]) = (0,0);
		(Bmult[24] => Cmult[29]) = (0,0);
		(Bmult[25] => Cmult[29]) = (0,0);
		(Bmult[26] => Cmult[29]) = (0,0);
		(Bmult[27] => Cmult[29]) = (0,0);
		(Bmult[28] => Cmult[29]) = (0,0);
		(Bmult[29] => Cmult[29]) = (0,0);
		(Bmult[30] => Cmult[29]) = (0,0);
		(Bmult[31] => Cmult[29]) = (0,0);		
		(Valid_mult[0] => Cmult[29]) = (0,0);
		(Valid_mult[1] => Cmult[29]) = (0,0);
		(sel_mul_32x32 => Cmult[29]) = (0,0);	
		(Amult[0]  => Cmult[30]) = (0,0);
		(Amult[1]  => Cmult[30]) = (0,0);
		(Amult[2]  => Cmult[30]) = (0,0);
		(Amult[3]  => Cmult[30]) = (0,0);
		(Amult[4]  => Cmult[30]) = (0,0);
		(Amult[5]  => Cmult[30]) = (0,0);
		(Amult[6]  => Cmult[30]) = (0,0);
		(Amult[7]  => Cmult[30]) = (0,0);
		(Amult[8]  => Cmult[30]) = (0,0);
		(Amult[9]  => Cmult[30]) = (0,0);
		(Amult[10] => Cmult[30]) = (0,0);
		(Amult[11] => Cmult[30]) = (0,0);
		(Amult[12] => Cmult[30]) = (0,0);
		(Amult[13] => Cmult[30]) = (0,0);
		(Amult[14] => Cmult[30]) = (0,0);
		(Amult[15] => Cmult[30]) = (0,0);
		(Amult[16] => Cmult[30]) = (0,0);
		(Amult[17] => Cmult[30]) = (0,0);
		(Amult[18] => Cmult[30]) = (0,0);
		(Amult[19] => Cmult[30]) = (0,0);
		(Amult[20] => Cmult[30]) = (0,0);
		(Amult[21] => Cmult[30]) = (0,0);
		(Amult[22] => Cmult[30]) = (0,0);
		(Amult[23] => Cmult[30]) = (0,0);
		(Amult[24] => Cmult[30]) = (0,0);
		(Amult[25] => Cmult[30]) = (0,0);
		(Amult[26] => Cmult[30]) = (0,0);
		(Amult[27] => Cmult[30]) = (0,0);
		(Amult[28] => Cmult[30]) = (0,0);
		(Amult[29] => Cmult[30]) = (0,0);
		(Amult[30] => Cmult[30]) = (0,0);
		(Amult[31] => Cmult[30]) = (0,0);
		(Bmult[0]  => Cmult[30]) = (0,0);
		(Bmult[1]  => Cmult[30]) = (0,0);
		(Bmult[2]  => Cmult[30]) = (0,0);
		(Bmult[3]  => Cmult[30]) = (0,0);
		(Bmult[4]  => Cmult[30]) = (0,0);
		(Bmult[5]  => Cmult[30]) = (0,0);
		(Bmult[6]  => Cmult[30]) = (0,0);
		(Bmult[7]  => Cmult[30]) = (0,0);
		(Bmult[8]  => Cmult[30]) = (0,0);
		(Bmult[9]  => Cmult[30]) = (0,0);
		(Bmult[10] => Cmult[30]) = (0,0);
		(Bmult[11] => Cmult[30]) = (0,0);
		(Bmult[12] => Cmult[30]) = (0,0);
		(Bmult[13] => Cmult[30]) = (0,0);
		(Bmult[14] => Cmult[30]) = (0,0);
		(Bmult[15] => Cmult[30]) = (0,0);
		(Bmult[16] => Cmult[30]) = (0,0);
		(Bmult[17] => Cmult[30]) = (0,0);
		(Bmult[18] => Cmult[30]) = (0,0);
		(Bmult[19] => Cmult[30]) = (0,0);
		(Bmult[20] => Cmult[30]) = (0,0);
		(Bmult[21] => Cmult[30]) = (0,0);
		(Bmult[22] => Cmult[30]) = (0,0);
		(Bmult[23] => Cmult[30]) = (0,0);
		(Bmult[24] => Cmult[30]) = (0,0);
		(Bmult[25] => Cmult[30]) = (0,0);
		(Bmult[26] => Cmult[30]) = (0,0);
		(Bmult[27] => Cmult[30]) = (0,0);
		(Bmult[28] => Cmult[30]) = (0,0);
		(Bmult[29] => Cmult[30]) = (0,0);
		(Bmult[30] => Cmult[30]) = (0,0);
		(Bmult[31] => Cmult[30]) = (0,0);		
		(Valid_mult[0] => Cmult[30]) = (0,0);
		(Valid_mult[1] => Cmult[30]) = (0,0);
		(sel_mul_32x32 => Cmult[30]) = (0,0);
		(Amult[0]  => Cmult[31]) = (0,0);
		(Amult[1]  => Cmult[31]) = (0,0);
		(Amult[2]  => Cmult[31]) = (0,0);
		(Amult[3]  => Cmult[31]) = (0,0);
		(Amult[4]  => Cmult[31]) = (0,0);
		(Amult[5]  => Cmult[31]) = (0,0);
		(Amult[6]  => Cmult[31]) = (0,0);
		(Amult[7]  => Cmult[31]) = (0,0);
		(Amult[8]  => Cmult[31]) = (0,0);
		(Amult[9]  => Cmult[31]) = (0,0);
		(Amult[10] => Cmult[31]) = (0,0);
		(Amult[11] => Cmult[31]) = (0,0);
		(Amult[12] => Cmult[31]) = (0,0);
		(Amult[13] => Cmult[31]) = (0,0);
		(Amult[14] => Cmult[31]) = (0,0);
		(Amult[15] => Cmult[31]) = (0,0);
		(Amult[16] => Cmult[31]) = (0,0);
		(Amult[17] => Cmult[31]) = (0,0);
		(Amult[18] => Cmult[31]) = (0,0);
		(Amult[19] => Cmult[31]) = (0,0);
		(Amult[20] => Cmult[31]) = (0,0);
		(Amult[21] => Cmult[31]) = (0,0);
		(Amult[22] => Cmult[31]) = (0,0);
		(Amult[23] => Cmult[31]) = (0,0);
		(Amult[24] => Cmult[31]) = (0,0);
		(Amult[25] => Cmult[31]) = (0,0);
		(Amult[26] => Cmult[31]) = (0,0);
		(Amult[27] => Cmult[31]) = (0,0);
		(Amult[28] => Cmult[31]) = (0,0);
		(Amult[29] => Cmult[31]) = (0,0);
		(Amult[30] => Cmult[31]) = (0,0);
		(Amult[31] => Cmult[31]) = (0,0);
		(Bmult[0]  => Cmult[31]) = (0,0);
		(Bmult[1]  => Cmult[31]) = (0,0);
		(Bmult[2]  => Cmult[31]) = (0,0);
		(Bmult[3]  => Cmult[31]) = (0,0);
		(Bmult[4]  => Cmult[31]) = (0,0);
		(Bmult[5]  => Cmult[31]) = (0,0);
		(Bmult[6]  => Cmult[31]) = (0,0);
		(Bmult[7]  => Cmult[31]) = (0,0);
		(Bmult[8]  => Cmult[31]) = (0,0);
		(Bmult[9]  => Cmult[31]) = (0,0);
		(Bmult[10] => Cmult[31]) = (0,0);
		(Bmult[11] => Cmult[31]) = (0,0);
		(Bmult[12] => Cmult[31]) = (0,0);
		(Bmult[13] => Cmult[31]) = (0,0);
		(Bmult[14] => Cmult[31]) = (0,0);
		(Bmult[15] => Cmult[31]) = (0,0);
		(Bmult[16] => Cmult[31]) = (0,0);
		(Bmult[17] => Cmult[31]) = (0,0);
		(Bmult[18] => Cmult[31]) = (0,0);
		(Bmult[19] => Cmult[31]) = (0,0);
		(Bmult[20] => Cmult[31]) = (0,0);
		(Bmult[21] => Cmult[31]) = (0,0);
		(Bmult[22] => Cmult[31]) = (0,0);
		(Bmult[23] => Cmult[31]) = (0,0);
		(Bmult[24] => Cmult[31]) = (0,0);
		(Bmult[25] => Cmult[31]) = (0,0);
		(Bmult[26] => Cmult[31]) = (0,0);
		(Bmult[27] => Cmult[31]) = (0,0);
		(Bmult[28] => Cmult[31]) = (0,0);
		(Bmult[29] => Cmult[31]) = (0,0);
		(Bmult[30] => Cmult[31]) = (0,0);
		(Bmult[31] => Cmult[31]) = (0,0);		
		(Valid_mult[0] => Cmult[31]) = (0,0);
		(Valid_mult[1] => Cmult[31]) = (0,0);
		(sel_mul_32x32 => Cmult[31]) = (0,0);
		(Amult[0]  => Cmult[32]) = (0,0);
		(Amult[1]  => Cmult[32]) = (0,0);
		(Amult[2]  => Cmult[32]) = (0,0);
		(Amult[3]  => Cmult[32]) = (0,0);
		(Amult[4]  => Cmult[32]) = (0,0);
		(Amult[5]  => Cmult[32]) = (0,0);
		(Amult[6]  => Cmult[32]) = (0,0);
		(Amult[7]  => Cmult[32]) = (0,0);
		(Amult[8]  => Cmult[32]) = (0,0);
		(Amult[9]  => Cmult[32]) = (0,0);
		(Amult[10] => Cmult[32]) = (0,0);
		(Amult[11] => Cmult[32]) = (0,0);
		(Amult[12] => Cmult[32]) = (0,0);
		(Amult[13] => Cmult[32]) = (0,0);
		(Amult[14] => Cmult[32]) = (0,0);
		(Amult[15] => Cmult[32]) = (0,0);
		(Amult[16] => Cmult[32]) = (0,0);
		(Amult[17] => Cmult[32]) = (0,0);
		(Amult[18] => Cmult[32]) = (0,0);
		(Amult[19] => Cmult[32]) = (0,0);
		(Amult[20] => Cmult[32]) = (0,0);
		(Amult[21] => Cmult[32]) = (0,0);
		(Amult[22] => Cmult[32]) = (0,0);
		(Amult[23] => Cmult[32]) = (0,0);
		(Amult[24] => Cmult[32]) = (0,0);
		(Amult[25] => Cmult[32]) = (0,0);
		(Amult[26] => Cmult[32]) = (0,0);
		(Amult[27] => Cmult[32]) = (0,0);
		(Amult[28] => Cmult[32]) = (0,0);
		(Amult[29] => Cmult[32]) = (0,0);
		(Amult[30] => Cmult[32]) = (0,0);
		(Amult[31] => Cmult[32]) = (0,0);
		(Bmult[0]  => Cmult[32]) = (0,0);
		(Bmult[1]  => Cmult[32]) = (0,0);
		(Bmult[2]  => Cmult[32]) = (0,0);
		(Bmult[3]  => Cmult[32]) = (0,0);
		(Bmult[4]  => Cmult[32]) = (0,0);
		(Bmult[5]  => Cmult[32]) = (0,0);
		(Bmult[6]  => Cmult[32]) = (0,0);
		(Bmult[7]  => Cmult[32]) = (0,0);
		(Bmult[8]  => Cmult[32]) = (0,0);
		(Bmult[9]  => Cmult[32]) = (0,0);
		(Bmult[10] => Cmult[32]) = (0,0);
		(Bmult[11] => Cmult[32]) = (0,0);
		(Bmult[12] => Cmult[32]) = (0,0);
		(Bmult[13] => Cmult[32]) = (0,0);
		(Bmult[14] => Cmult[32]) = (0,0);
		(Bmult[15] => Cmult[32]) = (0,0);
		(Bmult[16] => Cmult[32]) = (0,0);
		(Bmult[17] => Cmult[32]) = (0,0);
		(Bmult[18] => Cmult[32]) = (0,0);
		(Bmult[19] => Cmult[32]) = (0,0);
		(Bmult[20] => Cmult[32]) = (0,0);
		(Bmult[21] => Cmult[32]) = (0,0);
		(Bmult[22] => Cmult[32]) = (0,0);
		(Bmult[23] => Cmult[32]) = (0,0);
		(Bmult[24] => Cmult[32]) = (0,0);
		(Bmult[25] => Cmult[32]) = (0,0);
		(Bmult[26] => Cmult[32]) = (0,0);
		(Bmult[27] => Cmult[32]) = (0,0);
		(Bmult[28] => Cmult[32]) = (0,0);
		(Bmult[29] => Cmult[32]) = (0,0);
		(Bmult[30] => Cmult[32]) = (0,0);
		(Bmult[31] => Cmult[32]) = (0,0);		
		(Valid_mult[0] => Cmult[32]) = (0,0);
		(Valid_mult[1] => Cmult[32]) = (0,0);
		(sel_mul_32x32 => Cmult[32]) = (0,0);
		(Amult[0]  => Cmult[33]) = (0,0);
		(Amult[1]  => Cmult[33]) = (0,0);
		(Amult[2]  => Cmult[33]) = (0,0);
		(Amult[3]  => Cmult[33]) = (0,0);
		(Amult[4]  => Cmult[33]) = (0,0);
		(Amult[5]  => Cmult[33]) = (0,0);
		(Amult[6]  => Cmult[33]) = (0,0);
		(Amult[7]  => Cmult[33]) = (0,0);
		(Amult[8]  => Cmult[33]) = (0,0);
		(Amult[9]  => Cmult[33]) = (0,0);
		(Amult[10] => Cmult[33]) = (0,0);
		(Amult[11] => Cmult[33]) = (0,0);
		(Amult[12] => Cmult[33]) = (0,0);
		(Amult[13] => Cmult[33]) = (0,0);
		(Amult[14] => Cmult[33]) = (0,0);
		(Amult[15] => Cmult[33]) = (0,0);
		(Amult[16] => Cmult[33]) = (0,0);
		(Amult[17] => Cmult[33]) = (0,0);
		(Amult[18] => Cmult[33]) = (0,0);
		(Amult[19] => Cmult[33]) = (0,0);
		(Amult[20] => Cmult[33]) = (0,0);
		(Amult[21] => Cmult[33]) = (0,0);
		(Amult[22] => Cmult[33]) = (0,0);
		(Amult[23] => Cmult[33]) = (0,0);
		(Amult[24] => Cmult[33]) = (0,0);
		(Amult[25] => Cmult[33]) = (0,0);
		(Amult[26] => Cmult[33]) = (0,0);
		(Amult[27] => Cmult[33]) = (0,0);
		(Amult[28] => Cmult[33]) = (0,0);
		(Amult[29] => Cmult[33]) = (0,0);
		(Amult[30] => Cmult[33]) = (0,0);
		(Amult[31] => Cmult[33]) = (0,0);
		(Bmult[0]  => Cmult[33]) = (0,0);
		(Bmult[1]  => Cmult[33]) = (0,0);
		(Bmult[2]  => Cmult[33]) = (0,0);
		(Bmult[3]  => Cmult[33]) = (0,0);
		(Bmult[4]  => Cmult[33]) = (0,0);
		(Bmult[5]  => Cmult[33]) = (0,0);
		(Bmult[6]  => Cmult[33]) = (0,0);
		(Bmult[7]  => Cmult[33]) = (0,0);
		(Bmult[8]  => Cmult[33]) = (0,0);
		(Bmult[9]  => Cmult[33]) = (0,0);
		(Bmult[10] => Cmult[33]) = (0,0);
		(Bmult[11] => Cmult[33]) = (0,0);
		(Bmult[12] => Cmult[33]) = (0,0);
		(Bmult[13] => Cmult[33]) = (0,0);
		(Bmult[14] => Cmult[33]) = (0,0);
		(Bmult[15] => Cmult[33]) = (0,0);
		(Bmult[16] => Cmult[33]) = (0,0);
		(Bmult[17] => Cmult[33]) = (0,0);
		(Bmult[18] => Cmult[33]) = (0,0);
		(Bmult[19] => Cmult[33]) = (0,0);
		(Bmult[20] => Cmult[33]) = (0,0);
		(Bmult[21] => Cmult[33]) = (0,0);
		(Bmult[22] => Cmult[33]) = (0,0);
		(Bmult[23] => Cmult[33]) = (0,0);
		(Bmult[24] => Cmult[33]) = (0,0);
		(Bmult[25] => Cmult[33]) = (0,0);
		(Bmult[26] => Cmult[33]) = (0,0);
		(Bmult[27] => Cmult[33]) = (0,0);
		(Bmult[28] => Cmult[33]) = (0,0);
		(Bmult[29] => Cmult[33]) = (0,0);
		(Bmult[30] => Cmult[33]) = (0,0);
		(Bmult[31] => Cmult[33]) = (0,0);		
		(Valid_mult[0] => Cmult[33]) = (0,0);
		(Valid_mult[1] => Cmult[33]) = (0,0);
		(sel_mul_32x32 => Cmult[33]) = (0,0);
		(Amult[0]  => Cmult[34]) = (0,0);
		(Amult[1]  => Cmult[34]) = (0,0);
		(Amult[2]  => Cmult[34]) = (0,0);
		(Amult[3]  => Cmult[34]) = (0,0);
		(Amult[4]  => Cmult[34]) = (0,0);
		(Amult[5]  => Cmult[34]) = (0,0);
		(Amult[6]  => Cmult[34]) = (0,0);
		(Amult[7]  => Cmult[34]) = (0,0);
		(Amult[8]  => Cmult[34]) = (0,0);
		(Amult[9]  => Cmult[34]) = (0,0);
		(Amult[10] => Cmult[34]) = (0,0);
		(Amult[11] => Cmult[34]) = (0,0);
		(Amult[12] => Cmult[34]) = (0,0);
		(Amult[13] => Cmult[34]) = (0,0);
		(Amult[14] => Cmult[34]) = (0,0);
		(Amult[15] => Cmult[34]) = (0,0);
		(Amult[16] => Cmult[34]) = (0,0);
		(Amult[17] => Cmult[34]) = (0,0);
		(Amult[18] => Cmult[34]) = (0,0);
		(Amult[19] => Cmult[34]) = (0,0);
		(Amult[20] => Cmult[34]) = (0,0);
		(Amult[21] => Cmult[34]) = (0,0);
		(Amult[22] => Cmult[34]) = (0,0);
		(Amult[23] => Cmult[34]) = (0,0);
		(Amult[24] => Cmult[34]) = (0,0);
		(Amult[25] => Cmult[34]) = (0,0);
		(Amult[26] => Cmult[34]) = (0,0);
		(Amult[27] => Cmult[34]) = (0,0);
		(Amult[28] => Cmult[34]) = (0,0);
		(Amult[29] => Cmult[34]) = (0,0);
		(Amult[30] => Cmult[34]) = (0,0);
		(Amult[31] => Cmult[34]) = (0,0);
		(Bmult[0]  => Cmult[34]) = (0,0);
		(Bmult[1]  => Cmult[34]) = (0,0);
		(Bmult[2]  => Cmult[34]) = (0,0);
		(Bmult[3]  => Cmult[34]) = (0,0);
		(Bmult[4]  => Cmult[34]) = (0,0);
		(Bmult[5]  => Cmult[34]) = (0,0);
		(Bmult[6]  => Cmult[34]) = (0,0);
		(Bmult[7]  => Cmult[34]) = (0,0);
		(Bmult[8]  => Cmult[34]) = (0,0);
		(Bmult[9]  => Cmult[34]) = (0,0);
		(Bmult[10] => Cmult[34]) = (0,0);
		(Bmult[11] => Cmult[34]) = (0,0);
		(Bmult[12] => Cmult[34]) = (0,0);
		(Bmult[13] => Cmult[34]) = (0,0);
		(Bmult[14] => Cmult[34]) = (0,0);
		(Bmult[15] => Cmult[34]) = (0,0);
		(Bmult[16] => Cmult[34]) = (0,0);
		(Bmult[17] => Cmult[34]) = (0,0);
		(Bmult[18] => Cmult[34]) = (0,0);
		(Bmult[19] => Cmult[34]) = (0,0);
		(Bmult[20] => Cmult[34]) = (0,0);
		(Bmult[21] => Cmult[34]) = (0,0);
		(Bmult[22] => Cmult[34]) = (0,0);
		(Bmult[23] => Cmult[34]) = (0,0);
		(Bmult[24] => Cmult[34]) = (0,0);
		(Bmult[25] => Cmult[34]) = (0,0);
		(Bmult[26] => Cmult[34]) = (0,0);
		(Bmult[27] => Cmult[34]) = (0,0);
		(Bmult[28] => Cmult[34]) = (0,0);
		(Bmult[29] => Cmult[34]) = (0,0);
		(Bmult[30] => Cmult[34]) = (0,0);
		(Bmult[31] => Cmult[34]) = (0,0);		
		(Valid_mult[0] => Cmult[34]) = (0,0);
		(Valid_mult[1] => Cmult[34]) = (0,0);
		(sel_mul_32x32 => Cmult[34]) = (0,0);
		(Amult[0]  => Cmult[35]) = (0,0);
		(Amult[1]  => Cmult[35]) = (0,0);
		(Amult[2]  => Cmult[35]) = (0,0);
		(Amult[3]  => Cmult[35]) = (0,0);
		(Amult[4]  => Cmult[35]) = (0,0);
		(Amult[5]  => Cmult[35]) = (0,0);
		(Amult[6]  => Cmult[35]) = (0,0);
		(Amult[7]  => Cmult[35]) = (0,0);
		(Amult[8]  => Cmult[35]) = (0,0);
		(Amult[9]  => Cmult[35]) = (0,0);
		(Amult[10] => Cmult[35]) = (0,0);
		(Amult[11] => Cmult[35]) = (0,0);
		(Amult[12] => Cmult[35]) = (0,0);
		(Amult[13] => Cmult[35]) = (0,0);
		(Amult[14] => Cmult[35]) = (0,0);
		(Amult[15] => Cmult[35]) = (0,0);
		(Amult[16] => Cmult[35]) = (0,0);
		(Amult[17] => Cmult[35]) = (0,0);
		(Amult[18] => Cmult[35]) = (0,0);
		(Amult[19] => Cmult[35]) = (0,0);
		(Amult[20] => Cmult[35]) = (0,0);
		(Amult[21] => Cmult[35]) = (0,0);
		(Amult[22] => Cmult[35]) = (0,0);
		(Amult[23] => Cmult[35]) = (0,0);
		(Amult[24] => Cmult[35]) = (0,0);
		(Amult[25] => Cmult[35]) = (0,0);
		(Amult[26] => Cmult[35]) = (0,0);
		(Amult[27] => Cmult[35]) = (0,0);
		(Amult[28] => Cmult[35]) = (0,0);
		(Amult[29] => Cmult[35]) = (0,0);
		(Amult[30] => Cmult[35]) = (0,0);
		(Amult[31] => Cmult[35]) = (0,0);
		(Bmult[0]  => Cmult[35]) = (0,0);
		(Bmult[1]  => Cmult[35]) = (0,0);
		(Bmult[2]  => Cmult[35]) = (0,0);
		(Bmult[3]  => Cmult[35]) = (0,0);
		(Bmult[4]  => Cmult[35]) = (0,0);
		(Bmult[5]  => Cmult[35]) = (0,0);
		(Bmult[6]  => Cmult[35]) = (0,0);
		(Bmult[7]  => Cmult[35]) = (0,0);
		(Bmult[8]  => Cmult[35]) = (0,0);
		(Bmult[9]  => Cmult[35]) = (0,0);
		(Bmult[10] => Cmult[35]) = (0,0);
		(Bmult[11] => Cmult[35]) = (0,0);
		(Bmult[12] => Cmult[35]) = (0,0);
		(Bmult[13] => Cmult[35]) = (0,0);
		(Bmult[14] => Cmult[35]) = (0,0);
		(Bmult[15] => Cmult[35]) = (0,0);
		(Bmult[16] => Cmult[35]) = (0,0);
		(Bmult[17] => Cmult[35]) = (0,0);
		(Bmult[18] => Cmult[35]) = (0,0);
		(Bmult[19] => Cmult[35]) = (0,0);
		(Bmult[20] => Cmult[35]) = (0,0);
		(Bmult[21] => Cmult[35]) = (0,0);
		(Bmult[22] => Cmult[35]) = (0,0);
		(Bmult[23] => Cmult[35]) = (0,0);
		(Bmult[24] => Cmult[35]) = (0,0);
		(Bmult[25] => Cmult[35]) = (0,0);
		(Bmult[26] => Cmult[35]) = (0,0);
		(Bmult[27] => Cmult[35]) = (0,0);
		(Bmult[28] => Cmult[35]) = (0,0);
		(Bmult[29] => Cmult[35]) = (0,0);
		(Bmult[30] => Cmult[35]) = (0,0);
		(Bmult[31] => Cmult[35]) = (0,0);		
		(Valid_mult[0] => Cmult[35]) = (0,0);
		(Valid_mult[1] => Cmult[35]) = (0,0);
		(sel_mul_32x32 => Cmult[35]) = (0,0);
		(Amult[0]  => Cmult[36]) = (0,0);
		(Amult[1]  => Cmult[36]) = (0,0);
		(Amult[2]  => Cmult[36]) = (0,0);
		(Amult[3]  => Cmult[36]) = (0,0);
		(Amult[4]  => Cmult[36]) = (0,0);
		(Amult[5]  => Cmult[36]) = (0,0);
		(Amult[6]  => Cmult[36]) = (0,0);
		(Amult[7]  => Cmult[36]) = (0,0);
		(Amult[8]  => Cmult[36]) = (0,0);
		(Amult[9]  => Cmult[36]) = (0,0);
		(Amult[10] => Cmult[36]) = (0,0);
		(Amult[11] => Cmult[36]) = (0,0);
		(Amult[12] => Cmult[36]) = (0,0);
		(Amult[13] => Cmult[36]) = (0,0);
		(Amult[14] => Cmult[36]) = (0,0);
		(Amult[15] => Cmult[36]) = (0,0);
		(Amult[16] => Cmult[36]) = (0,0);
		(Amult[17] => Cmult[36]) = (0,0);
		(Amult[18] => Cmult[36]) = (0,0);
		(Amult[19] => Cmult[36]) = (0,0);
		(Amult[20] => Cmult[36]) = (0,0);
		(Amult[21] => Cmult[36]) = (0,0);
		(Amult[22] => Cmult[36]) = (0,0);
		(Amult[23] => Cmult[36]) = (0,0);
		(Amult[24] => Cmult[36]) = (0,0);
		(Amult[25] => Cmult[36]) = (0,0);
		(Amult[26] => Cmult[36]) = (0,0);
		(Amult[27] => Cmult[36]) = (0,0);
		(Amult[28] => Cmult[36]) = (0,0);
		(Amult[29] => Cmult[36]) = (0,0);
		(Amult[30] => Cmult[36]) = (0,0);
		(Amult[31] => Cmult[36]) = (0,0);
		(Bmult[0]  => Cmult[36]) = (0,0);
		(Bmult[1]  => Cmult[36]) = (0,0);
		(Bmult[2]  => Cmult[36]) = (0,0);
		(Bmult[3]  => Cmult[36]) = (0,0);
		(Bmult[4]  => Cmult[36]) = (0,0);
		(Bmult[5]  => Cmult[36]) = (0,0);
		(Bmult[6]  => Cmult[36]) = (0,0);
		(Bmult[7]  => Cmult[36]) = (0,0);
		(Bmult[8]  => Cmult[36]) = (0,0);
		(Bmult[9]  => Cmult[36]) = (0,0);
		(Bmult[10] => Cmult[36]) = (0,0);
		(Bmult[11] => Cmult[36]) = (0,0);
		(Bmult[12] => Cmult[36]) = (0,0);
		(Bmult[13] => Cmult[36]) = (0,0);
		(Bmult[14] => Cmult[36]) = (0,0);
		(Bmult[15] => Cmult[36]) = (0,0);
		(Bmult[16] => Cmult[36]) = (0,0);
		(Bmult[17] => Cmult[36]) = (0,0);
		(Bmult[18] => Cmult[36]) = (0,0);
		(Bmult[19] => Cmult[36]) = (0,0);
		(Bmult[20] => Cmult[36]) = (0,0);
		(Bmult[21] => Cmult[36]) = (0,0);
		(Bmult[22] => Cmult[36]) = (0,0);
		(Bmult[23] => Cmult[36]) = (0,0);
		(Bmult[24] => Cmult[36]) = (0,0);
		(Bmult[25] => Cmult[36]) = (0,0);
		(Bmult[26] => Cmult[36]) = (0,0);
		(Bmult[27] => Cmult[36]) = (0,0);
		(Bmult[28] => Cmult[36]) = (0,0);
		(Bmult[29] => Cmult[36]) = (0,0);
		(Bmult[30] => Cmult[36]) = (0,0);
		(Bmult[31] => Cmult[36]) = (0,0);		
		(Valid_mult[0] => Cmult[36]) = (0,0);
		(Valid_mult[1] => Cmult[36]) = (0,0);
		(sel_mul_32x32 => Cmult[36]) = (0,0);
		(Amult[0]  => Cmult[37]) = (0,0);
		(Amult[1]  => Cmult[37]) = (0,0);
		(Amult[2]  => Cmult[37]) = (0,0);
		(Amult[3]  => Cmult[37]) = (0,0);
		(Amult[4]  => Cmult[37]) = (0,0);
		(Amult[5]  => Cmult[37]) = (0,0);
		(Amult[6]  => Cmult[37]) = (0,0);
		(Amult[7]  => Cmult[37]) = (0,0);
		(Amult[8]  => Cmult[37]) = (0,0);
		(Amult[9]  => Cmult[37]) = (0,0);
		(Amult[10] => Cmult[37]) = (0,0);
		(Amult[11] => Cmult[37]) = (0,0);
		(Amult[12] => Cmult[37]) = (0,0);
		(Amult[13] => Cmult[37]) = (0,0);
		(Amult[14] => Cmult[37]) = (0,0);
		(Amult[15] => Cmult[37]) = (0,0);
		(Amult[16] => Cmult[37]) = (0,0);
		(Amult[17] => Cmult[37]) = (0,0);
		(Amult[18] => Cmult[37]) = (0,0);
		(Amult[19] => Cmult[37]) = (0,0);
		(Amult[20] => Cmult[37]) = (0,0);
		(Amult[21] => Cmult[37]) = (0,0);
		(Amult[22] => Cmult[37]) = (0,0);
		(Amult[23] => Cmult[37]) = (0,0);
		(Amult[24] => Cmult[37]) = (0,0);
		(Amult[25] => Cmult[37]) = (0,0);
		(Amult[26] => Cmult[37]) = (0,0);
		(Amult[27] => Cmult[37]) = (0,0);
		(Amult[28] => Cmult[37]) = (0,0);
		(Amult[29] => Cmult[37]) = (0,0);
		(Amult[30] => Cmult[37]) = (0,0);
		(Amult[31] => Cmult[37]) = (0,0);
		(Bmult[0]  => Cmult[37]) = (0,0);
		(Bmult[1]  => Cmult[37]) = (0,0);
		(Bmult[2]  => Cmult[37]) = (0,0);
		(Bmult[3]  => Cmult[37]) = (0,0);
		(Bmult[4]  => Cmult[37]) = (0,0);
		(Bmult[5]  => Cmult[37]) = (0,0);
		(Bmult[6]  => Cmult[37]) = (0,0);
		(Bmult[7]  => Cmult[37]) = (0,0);
		(Bmult[8]  => Cmult[37]) = (0,0);
		(Bmult[9]  => Cmult[37]) = (0,0);
		(Bmult[10] => Cmult[37]) = (0,0);
		(Bmult[11] => Cmult[37]) = (0,0);
		(Bmult[12] => Cmult[37]) = (0,0);
		(Bmult[13] => Cmult[37]) = (0,0);
		(Bmult[14] => Cmult[37]) = (0,0);
		(Bmult[15] => Cmult[37]) = (0,0);
		(Bmult[16] => Cmult[37]) = (0,0);
		(Bmult[17] => Cmult[37]) = (0,0);
		(Bmult[18] => Cmult[37]) = (0,0);
		(Bmult[19] => Cmult[37]) = (0,0);
		(Bmult[20] => Cmult[37]) = (0,0);
		(Bmult[21] => Cmult[37]) = (0,0);
		(Bmult[22] => Cmult[37]) = (0,0);
		(Bmult[23] => Cmult[37]) = (0,0);
		(Bmult[24] => Cmult[37]) = (0,0);
		(Bmult[25] => Cmult[37]) = (0,0);
		(Bmult[26] => Cmult[37]) = (0,0);
		(Bmult[27] => Cmult[37]) = (0,0);
		(Bmult[28] => Cmult[37]) = (0,0);
		(Bmult[29] => Cmult[37]) = (0,0);
		(Bmult[30] => Cmult[37]) = (0,0);
		(Bmult[31] => Cmult[37]) = (0,0);		
		(Valid_mult[0] => Cmult[37]) = (0,0);
		(Valid_mult[1] => Cmult[37]) = (0,0);
		(sel_mul_32x32 => Cmult[37]) = (0,0);
		(Amult[0]  => Cmult[38]) = (0,0);
		(Amult[1]  => Cmult[38]) = (0,0);
		(Amult[2]  => Cmult[38]) = (0,0);
		(Amult[3]  => Cmult[38]) = (0,0);
		(Amult[4]  => Cmult[38]) = (0,0);
		(Amult[5]  => Cmult[38]) = (0,0);
		(Amult[6]  => Cmult[38]) = (0,0);
		(Amult[7]  => Cmult[38]) = (0,0);
		(Amult[8]  => Cmult[38]) = (0,0);
		(Amult[9]  => Cmult[38]) = (0,0);
		(Amult[10] => Cmult[38]) = (0,0);
		(Amult[11] => Cmult[38]) = (0,0);
		(Amult[12] => Cmult[38]) = (0,0);
		(Amult[13] => Cmult[38]) = (0,0);
		(Amult[14] => Cmult[38]) = (0,0);
		(Amult[15] => Cmult[38]) = (0,0);
		(Amult[16] => Cmult[38]) = (0,0);
		(Amult[17] => Cmult[38]) = (0,0);
		(Amult[18] => Cmult[38]) = (0,0);
		(Amult[19] => Cmult[38]) = (0,0);
		(Amult[20] => Cmult[38]) = (0,0);
		(Amult[21] => Cmult[38]) = (0,0);
		(Amult[22] => Cmult[38]) = (0,0);
		(Amult[23] => Cmult[38]) = (0,0);
		(Amult[24] => Cmult[38]) = (0,0);
		(Amult[25] => Cmult[38]) = (0,0);
		(Amult[26] => Cmult[38]) = (0,0);
		(Amult[27] => Cmult[38]) = (0,0);
		(Amult[28] => Cmult[38]) = (0,0);
		(Amult[29] => Cmult[38]) = (0,0);
		(Amult[30] => Cmult[38]) = (0,0);
		(Amult[31] => Cmult[38]) = (0,0);
		(Bmult[0]  => Cmult[38]) = (0,0);
		(Bmult[1]  => Cmult[38]) = (0,0);
		(Bmult[2]  => Cmult[38]) = (0,0);
		(Bmult[3]  => Cmult[38]) = (0,0);
		(Bmult[4]  => Cmult[38]) = (0,0);
		(Bmult[5]  => Cmult[38]) = (0,0);
		(Bmult[6]  => Cmult[38]) = (0,0);
		(Bmult[7]  => Cmult[38]) = (0,0);
		(Bmult[8]  => Cmult[38]) = (0,0);
		(Bmult[9]  => Cmult[38]) = (0,0);
		(Bmult[10] => Cmult[38]) = (0,0);
		(Bmult[11] => Cmult[38]) = (0,0);
		(Bmult[12] => Cmult[38]) = (0,0);
		(Bmult[13] => Cmult[38]) = (0,0);
		(Bmult[14] => Cmult[38]) = (0,0);
		(Bmult[15] => Cmult[38]) = (0,0);
		(Bmult[16] => Cmult[38]) = (0,0);
		(Bmult[17] => Cmult[38]) = (0,0);
		(Bmult[18] => Cmult[38]) = (0,0);
		(Bmult[19] => Cmult[38]) = (0,0);
		(Bmult[20] => Cmult[38]) = (0,0);
		(Bmult[21] => Cmult[38]) = (0,0);
		(Bmult[22] => Cmult[38]) = (0,0);
		(Bmult[23] => Cmult[38]) = (0,0);
		(Bmult[24] => Cmult[38]) = (0,0);
		(Bmult[25] => Cmult[38]) = (0,0);
		(Bmult[26] => Cmult[38]) = (0,0);
		(Bmult[27] => Cmult[38]) = (0,0);
		(Bmult[28] => Cmult[38]) = (0,0);
		(Bmult[29] => Cmult[38]) = (0,0);
		(Bmult[30] => Cmult[38]) = (0,0);
		(Bmult[31] => Cmult[38]) = (0,0);		
		(Valid_mult[0] => Cmult[38]) = (0,0);
		(Valid_mult[1] => Cmult[38]) = (0,0);
		(sel_mul_32x32 => Cmult[38]) = (0,0);	
		(Amult[0]  => Cmult[39]) = (0,0);
		(Amult[1]  => Cmult[39]) = (0,0);
		(Amult[2]  => Cmult[39]) = (0,0);
		(Amult[3]  => Cmult[39]) = (0,0);
		(Amult[4]  => Cmult[39]) = (0,0);
		(Amult[5]  => Cmult[39]) = (0,0);
		(Amult[6]  => Cmult[39]) = (0,0);
		(Amult[7]  => Cmult[39]) = (0,0);
		(Amult[8]  => Cmult[39]) = (0,0);
		(Amult[9]  => Cmult[39]) = (0,0);
		(Amult[10] => Cmult[39]) = (0,0);
		(Amult[11] => Cmult[39]) = (0,0);
		(Amult[12] => Cmult[39]) = (0,0);
		(Amult[13] => Cmult[39]) = (0,0);
		(Amult[14] => Cmult[39]) = (0,0);
		(Amult[15] => Cmult[39]) = (0,0);
		(Amult[16] => Cmult[39]) = (0,0);
		(Amult[17] => Cmult[39]) = (0,0);
		(Amult[18] => Cmult[39]) = (0,0);
		(Amult[19] => Cmult[39]) = (0,0);
		(Amult[20] => Cmult[39]) = (0,0);
		(Amult[21] => Cmult[39]) = (0,0);
		(Amult[22] => Cmult[39]) = (0,0);
		(Amult[23] => Cmult[39]) = (0,0);
		(Amult[24] => Cmult[39]) = (0,0);
		(Amult[25] => Cmult[39]) = (0,0);
		(Amult[26] => Cmult[39]) = (0,0);
		(Amult[27] => Cmult[39]) = (0,0);
		(Amult[28] => Cmult[39]) = (0,0);
		(Amult[29] => Cmult[39]) = (0,0);
		(Amult[30] => Cmult[39]) = (0,0);
		(Amult[31] => Cmult[39]) = (0,0);
		(Bmult[0]  => Cmult[39]) = (0,0);
		(Bmult[1]  => Cmult[39]) = (0,0);
		(Bmult[2]  => Cmult[39]) = (0,0);
		(Bmult[3]  => Cmult[39]) = (0,0);
		(Bmult[4]  => Cmult[39]) = (0,0);
		(Bmult[5]  => Cmult[39]) = (0,0);
		(Bmult[6]  => Cmult[39]) = (0,0);
		(Bmult[7]  => Cmult[39]) = (0,0);
		(Bmult[8]  => Cmult[39]) = (0,0);
		(Bmult[9]  => Cmult[39]) = (0,0);
		(Bmult[10] => Cmult[39]) = (0,0);
		(Bmult[11] => Cmult[39]) = (0,0);
		(Bmult[12] => Cmult[39]) = (0,0);
		(Bmult[13] => Cmult[39]) = (0,0);
		(Bmult[14] => Cmult[39]) = (0,0);
		(Bmult[15] => Cmult[39]) = (0,0);
		(Bmult[16] => Cmult[39]) = (0,0);
		(Bmult[17] => Cmult[39]) = (0,0);
		(Bmult[18] => Cmult[39]) = (0,0);
		(Bmult[19] => Cmult[39]) = (0,0);
		(Bmult[20] => Cmult[39]) = (0,0);
		(Bmult[21] => Cmult[39]) = (0,0);
		(Bmult[22] => Cmult[39]) = (0,0);
		(Bmult[23] => Cmult[39]) = (0,0);
		(Bmult[24] => Cmult[39]) = (0,0);
		(Bmult[25] => Cmult[39]) = (0,0);
		(Bmult[26] => Cmult[39]) = (0,0);
		(Bmult[27] => Cmult[39]) = (0,0);
		(Bmult[28] => Cmult[39]) = (0,0);
		(Bmult[29] => Cmult[39]) = (0,0);
		(Bmult[30] => Cmult[39]) = (0,0);
		(Bmult[31] => Cmult[39]) = (0,0);		
		(Valid_mult[0] => Cmult[39]) = (0,0);
		(Valid_mult[1] => Cmult[39]) = (0,0);
		(sel_mul_32x32 => Cmult[39]) = (0,0);
		(Amult[0]  => Cmult[40]) = (0,0);
		(Amult[1]  => Cmult[40]) = (0,0);
		(Amult[2]  => Cmult[40]) = (0,0);
		(Amult[3]  => Cmult[40]) = (0,0);
		(Amult[4]  => Cmult[40]) = (0,0);
		(Amult[5]  => Cmult[40]) = (0,0);
		(Amult[6]  => Cmult[40]) = (0,0);
		(Amult[7]  => Cmult[40]) = (0,0);
		(Amult[8]  => Cmult[40]) = (0,0);
		(Amult[9]  => Cmult[40]) = (0,0);
		(Amult[10] => Cmult[40]) = (0,0);
		(Amult[11] => Cmult[40]) = (0,0);
		(Amult[12] => Cmult[40]) = (0,0);
		(Amult[13] => Cmult[40]) = (0,0);
		(Amult[14] => Cmult[40]) = (0,0);
		(Amult[15] => Cmult[40]) = (0,0);
		(Amult[16] => Cmult[40]) = (0,0);
		(Amult[17] => Cmult[40]) = (0,0);
		(Amult[18] => Cmult[40]) = (0,0);
		(Amult[19] => Cmult[40]) = (0,0);
		(Amult[20] => Cmult[40]) = (0,0);
		(Amult[21] => Cmult[40]) = (0,0);
		(Amult[22] => Cmult[40]) = (0,0);
		(Amult[23] => Cmult[40]) = (0,0);
		(Amult[24] => Cmult[40]) = (0,0);
		(Amult[25] => Cmult[40]) = (0,0);
		(Amult[26] => Cmult[40]) = (0,0);
		(Amult[27] => Cmult[40]) = (0,0);
		(Amult[28] => Cmult[40]) = (0,0);
		(Amult[29] => Cmult[40]) = (0,0);
		(Amult[30] => Cmult[40]) = (0,0);
		(Amult[31] => Cmult[40]) = (0,0);
		(Bmult[0]  => Cmult[40]) = (0,0);
		(Bmult[1]  => Cmult[40]) = (0,0);
		(Bmult[2]  => Cmult[40]) = (0,0);
		(Bmult[3]  => Cmult[40]) = (0,0);
		(Bmult[4]  => Cmult[40]) = (0,0);
		(Bmult[5]  => Cmult[40]) = (0,0);
		(Bmult[6]  => Cmult[40]) = (0,0);
		(Bmult[7]  => Cmult[40]) = (0,0);
		(Bmult[8]  => Cmult[40]) = (0,0);
		(Bmult[9]  => Cmult[40]) = (0,0);
		(Bmult[10] => Cmult[40]) = (0,0);
		(Bmult[11] => Cmult[40]) = (0,0);
		(Bmult[12] => Cmult[40]) = (0,0);
		(Bmult[13] => Cmult[40]) = (0,0);
		(Bmult[14] => Cmult[40]) = (0,0);
		(Bmult[15] => Cmult[40]) = (0,0);
		(Bmult[16] => Cmult[40]) = (0,0);
		(Bmult[17] => Cmult[40]) = (0,0);
		(Bmult[18] => Cmult[40]) = (0,0);
		(Bmult[19] => Cmult[40]) = (0,0);
		(Bmult[20] => Cmult[40]) = (0,0);
		(Bmult[21] => Cmult[40]) = (0,0);
		(Bmult[22] => Cmult[40]) = (0,0);
		(Bmult[23] => Cmult[40]) = (0,0);
		(Bmult[24] => Cmult[40]) = (0,0);
		(Bmult[25] => Cmult[40]) = (0,0);
		(Bmult[26] => Cmult[40]) = (0,0);
		(Bmult[27] => Cmult[40]) = (0,0);
		(Bmult[28] => Cmult[40]) = (0,0);
		(Bmult[29] => Cmult[40]) = (0,0);
		(Bmult[30] => Cmult[40]) = (0,0);
		(Bmult[31] => Cmult[40]) = (0,0);		
		(Valid_mult[0] => Cmult[40]) = (0,0);
		(Valid_mult[1] => Cmult[40]) = (0,0);
		(sel_mul_32x32 => Cmult[40]) = (0,0);
		(Amult[0]  => Cmult[41]) = (0,0);
		(Amult[1]  => Cmult[41]) = (0,0);
		(Amult[2]  => Cmult[41]) = (0,0);
		(Amult[3]  => Cmult[41]) = (0,0);
		(Amult[4]  => Cmult[41]) = (0,0);
		(Amult[5]  => Cmult[41]) = (0,0);
		(Amult[6]  => Cmult[41]) = (0,0);
		(Amult[7]  => Cmult[41]) = (0,0);
		(Amult[8]  => Cmult[41]) = (0,0);
		(Amult[9]  => Cmult[41]) = (0,0);
		(Amult[10] => Cmult[41]) = (0,0);
		(Amult[11] => Cmult[41]) = (0,0);
		(Amult[12] => Cmult[41]) = (0,0);
		(Amult[13] => Cmult[41]) = (0,0);
		(Amult[14] => Cmult[41]) = (0,0);
		(Amult[15] => Cmult[41]) = (0,0);
		(Amult[16] => Cmult[41]) = (0,0);
		(Amult[17] => Cmult[41]) = (0,0);
		(Amult[18] => Cmult[41]) = (0,0);
		(Amult[19] => Cmult[41]) = (0,0);
		(Amult[20] => Cmult[41]) = (0,0);
		(Amult[21] => Cmult[41]) = (0,0);
		(Amult[22] => Cmult[41]) = (0,0);
		(Amult[23] => Cmult[41]) = (0,0);
		(Amult[24] => Cmult[41]) = (0,0);
		(Amult[25] => Cmult[41]) = (0,0);
		(Amult[26] => Cmult[41]) = (0,0);
		(Amult[27] => Cmult[41]) = (0,0);
		(Amult[28] => Cmult[41]) = (0,0);
		(Amult[29] => Cmult[41]) = (0,0);
		(Amult[30] => Cmult[41]) = (0,0);
		(Amult[31] => Cmult[41]) = (0,0);
		(Bmult[0]  => Cmult[41]) = (0,0);
		(Bmult[1]  => Cmult[41]) = (0,0);
		(Bmult[2]  => Cmult[41]) = (0,0);
		(Bmult[3]  => Cmult[41]) = (0,0);
		(Bmult[4]  => Cmult[41]) = (0,0);
		(Bmult[5]  => Cmult[41]) = (0,0);
		(Bmult[6]  => Cmult[41]) = (0,0);
		(Bmult[7]  => Cmult[41]) = (0,0);
		(Bmult[8]  => Cmult[41]) = (0,0);
		(Bmult[9]  => Cmult[41]) = (0,0);
		(Bmult[10] => Cmult[41]) = (0,0);
		(Bmult[11] => Cmult[41]) = (0,0);
		(Bmult[12] => Cmult[41]) = (0,0);
		(Bmult[13] => Cmult[41]) = (0,0);
		(Bmult[14] => Cmult[41]) = (0,0);
		(Bmult[15] => Cmult[41]) = (0,0);
		(Bmult[16] => Cmult[41]) = (0,0);
		(Bmult[17] => Cmult[41]) = (0,0);
		(Bmult[18] => Cmult[41]) = (0,0);
		(Bmult[19] => Cmult[41]) = (0,0);
		(Bmult[20] => Cmult[41]) = (0,0);
		(Bmult[21] => Cmult[41]) = (0,0);
		(Bmult[22] => Cmult[41]) = (0,0);
		(Bmult[23] => Cmult[41]) = (0,0);
		(Bmult[24] => Cmult[41]) = (0,0);
		(Bmult[25] => Cmult[41]) = (0,0);
		(Bmult[26] => Cmult[41]) = (0,0);
		(Bmult[27] => Cmult[41]) = (0,0);
		(Bmult[28] => Cmult[41]) = (0,0);
		(Bmult[29] => Cmult[41]) = (0,0);
		(Bmult[30] => Cmult[41]) = (0,0);
		(Bmult[31] => Cmult[41]) = (0,0);		
		(Valid_mult[0] => Cmult[41]) = (0,0);
		(Valid_mult[1] => Cmult[41]) = (0,0);
		(sel_mul_32x32 => Cmult[41]) = (0,0);
		(Amult[0]  => Cmult[42]) = (0,0);
		(Amult[1]  => Cmult[42]) = (0,0);
		(Amult[2]  => Cmult[42]) = (0,0);
		(Amult[3]  => Cmult[42]) = (0,0);
		(Amult[4]  => Cmult[42]) = (0,0);
		(Amult[5]  => Cmult[42]) = (0,0);
		(Amult[6]  => Cmult[42]) = (0,0);
		(Amult[7]  => Cmult[42]) = (0,0);
		(Amult[8]  => Cmult[42]) = (0,0);
		(Amult[9]  => Cmult[42]) = (0,0);
		(Amult[10] => Cmult[42]) = (0,0);
		(Amult[11] => Cmult[42]) = (0,0);
		(Amult[12] => Cmult[42]) = (0,0);
		(Amult[13] => Cmult[42]) = (0,0);
		(Amult[14] => Cmult[42]) = (0,0);
		(Amult[15] => Cmult[42]) = (0,0);
		(Amult[16] => Cmult[42]) = (0,0);
		(Amult[17] => Cmult[42]) = (0,0);
		(Amult[18] => Cmult[42]) = (0,0);
		(Amult[19] => Cmult[42]) = (0,0);
		(Amult[20] => Cmult[42]) = (0,0);
		(Amult[21] => Cmult[42]) = (0,0);
		(Amult[22] => Cmult[42]) = (0,0);
		(Amult[23] => Cmult[42]) = (0,0);
		(Amult[24] => Cmult[42]) = (0,0);
		(Amult[25] => Cmult[42]) = (0,0);
		(Amult[26] => Cmult[42]) = (0,0);
		(Amult[27] => Cmult[42]) = (0,0);
		(Amult[28] => Cmult[42]) = (0,0);
		(Amult[29] => Cmult[42]) = (0,0);
		(Amult[30] => Cmult[42]) = (0,0);
		(Amult[31] => Cmult[42]) = (0,0);
		(Bmult[0]  => Cmult[42]) = (0,0);
		(Bmult[1]  => Cmult[42]) = (0,0);
		(Bmult[2]  => Cmult[42]) = (0,0);
		(Bmult[3]  => Cmult[42]) = (0,0);
		(Bmult[4]  => Cmult[42]) = (0,0);
		(Bmult[5]  => Cmult[42]) = (0,0);
		(Bmult[6]  => Cmult[42]) = (0,0);
		(Bmult[7]  => Cmult[42]) = (0,0);
		(Bmult[8]  => Cmult[42]) = (0,0);
		(Bmult[9]  => Cmult[42]) = (0,0);
		(Bmult[10] => Cmult[42]) = (0,0);
		(Bmult[11] => Cmult[42]) = (0,0);
		(Bmult[12] => Cmult[42]) = (0,0);
		(Bmult[13] => Cmult[42]) = (0,0);
		(Bmult[14] => Cmult[42]) = (0,0);
		(Bmult[15] => Cmult[42]) = (0,0);
		(Bmult[16] => Cmult[42]) = (0,0);
		(Bmult[17] => Cmult[42]) = (0,0);
		(Bmult[18] => Cmult[42]) = (0,0);
		(Bmult[19] => Cmult[42]) = (0,0);
		(Bmult[20] => Cmult[42]) = (0,0);
		(Bmult[21] => Cmult[42]) = (0,0);
		(Bmult[22] => Cmult[42]) = (0,0);
		(Bmult[23] => Cmult[42]) = (0,0);
		(Bmult[24] => Cmult[42]) = (0,0);
		(Bmult[25] => Cmult[42]) = (0,0);
		(Bmult[26] => Cmult[42]) = (0,0);
		(Bmult[27] => Cmult[42]) = (0,0);
		(Bmult[28] => Cmult[42]) = (0,0);
		(Bmult[29] => Cmult[42]) = (0,0);
		(Bmult[30] => Cmult[42]) = (0,0);
		(Bmult[31] => Cmult[42]) = (0,0);		
		(Valid_mult[0] => Cmult[42]) = (0,0);
		(Valid_mult[1] => Cmult[42]) = (0,0);
		(sel_mul_32x32 => Cmult[42]) = (0,0);
		(Amult[0]  => Cmult[43]) = (0,0);
		(Amult[1]  => Cmult[43]) = (0,0);
		(Amult[2]  => Cmult[43]) = (0,0);
		(Amult[3]  => Cmult[43]) = (0,0);
		(Amult[4]  => Cmult[43]) = (0,0);
		(Amult[5]  => Cmult[43]) = (0,0);
		(Amult[6]  => Cmult[43]) = (0,0);
		(Amult[7]  => Cmult[43]) = (0,0);
		(Amult[8]  => Cmult[43]) = (0,0);
		(Amult[9]  => Cmult[43]) = (0,0);
		(Amult[10] => Cmult[43]) = (0,0);
		(Amult[11] => Cmult[43]) = (0,0);
		(Amult[12] => Cmult[43]) = (0,0);
		(Amult[13] => Cmult[43]) = (0,0);
		(Amult[14] => Cmult[43]) = (0,0);
		(Amult[15] => Cmult[43]) = (0,0);
		(Amult[16] => Cmult[43]) = (0,0);
		(Amult[17] => Cmult[43]) = (0,0);
		(Amult[18] => Cmult[43]) = (0,0);
		(Amult[19] => Cmult[43]) = (0,0);
		(Amult[20] => Cmult[43]) = (0,0);
		(Amult[21] => Cmult[43]) = (0,0);
		(Amult[22] => Cmult[43]) = (0,0);
		(Amult[23] => Cmult[43]) = (0,0);
		(Amult[24] => Cmult[43]) = (0,0);
		(Amult[25] => Cmult[43]) = (0,0);
		(Amult[26] => Cmult[43]) = (0,0);
		(Amult[27] => Cmult[43]) = (0,0);
		(Amult[28] => Cmult[43]) = (0,0);
		(Amult[29] => Cmult[43]) = (0,0);
		(Amult[30] => Cmult[43]) = (0,0);
		(Amult[31] => Cmult[43]) = (0,0);
		(Bmult[0]  => Cmult[43]) = (0,0);
		(Bmult[1]  => Cmult[43]) = (0,0);
		(Bmult[2]  => Cmult[43]) = (0,0);
		(Bmult[3]  => Cmult[43]) = (0,0);
		(Bmult[4]  => Cmult[43]) = (0,0);
		(Bmult[5]  => Cmult[43]) = (0,0);
		(Bmult[6]  => Cmult[43]) = (0,0);
		(Bmult[7]  => Cmult[43]) = (0,0);
		(Bmult[8]  => Cmult[43]) = (0,0);
		(Bmult[9]  => Cmult[43]) = (0,0);
		(Bmult[10] => Cmult[43]) = (0,0);
		(Bmult[11] => Cmult[43]) = (0,0);
		(Bmult[12] => Cmult[43]) = (0,0);
		(Bmult[13] => Cmult[43]) = (0,0);
		(Bmult[14] => Cmult[43]) = (0,0);
		(Bmult[15] => Cmult[43]) = (0,0);
		(Bmult[16] => Cmult[43]) = (0,0);
		(Bmult[17] => Cmult[43]) = (0,0);
		(Bmult[18] => Cmult[43]) = (0,0);
		(Bmult[19] => Cmult[43]) = (0,0);
		(Bmult[20] => Cmult[43]) = (0,0);
		(Bmult[21] => Cmult[43]) = (0,0);
		(Bmult[22] => Cmult[43]) = (0,0);
		(Bmult[23] => Cmult[43]) = (0,0);
		(Bmult[24] => Cmult[43]) = (0,0);
		(Bmult[25] => Cmult[43]) = (0,0);
		(Bmult[26] => Cmult[43]) = (0,0);
		(Bmult[27] => Cmult[43]) = (0,0);
		(Bmult[28] => Cmult[43]) = (0,0);
		(Bmult[29] => Cmult[43]) = (0,0);
		(Bmult[30] => Cmult[43]) = (0,0);
		(Bmult[31] => Cmult[43]) = (0,0);		
		(Valid_mult[0] => Cmult[43]) = (0,0);
		(Valid_mult[1] => Cmult[43]) = (0,0);
		(sel_mul_32x32 => Cmult[43]) = (0,0);
		(Amult[0]  => Cmult[44]) = (0,0);
		(Amult[1]  => Cmult[44]) = (0,0);
		(Amult[2]  => Cmult[44]) = (0,0);
		(Amult[3]  => Cmult[44]) = (0,0);
		(Amult[4]  => Cmult[44]) = (0,0);
		(Amult[5]  => Cmult[44]) = (0,0);
		(Amult[6]  => Cmult[44]) = (0,0);
		(Amult[7]  => Cmult[44]) = (0,0);
		(Amult[8]  => Cmult[44]) = (0,0);
		(Amult[9]  => Cmult[44]) = (0,0);
		(Amult[10] => Cmult[44]) = (0,0);
		(Amult[11] => Cmult[44]) = (0,0);
		(Amult[12] => Cmult[44]) = (0,0);
		(Amult[13] => Cmult[44]) = (0,0);
		(Amult[14] => Cmult[44]) = (0,0);
		(Amult[15] => Cmult[44]) = (0,0);
		(Amult[16] => Cmult[44]) = (0,0);
		(Amult[17] => Cmult[44]) = (0,0);
		(Amult[18] => Cmult[44]) = (0,0);
		(Amult[19] => Cmult[44]) = (0,0);
		(Amult[20] => Cmult[44]) = (0,0);
		(Amult[21] => Cmult[44]) = (0,0);
		(Amult[22] => Cmult[44]) = (0,0);
		(Amult[23] => Cmult[44]) = (0,0);
		(Amult[24] => Cmult[44]) = (0,0);
		(Amult[25] => Cmult[44]) = (0,0);
		(Amult[26] => Cmult[44]) = (0,0);
		(Amult[27] => Cmult[44]) = (0,0);
		(Amult[28] => Cmult[44]) = (0,0);
		(Amult[29] => Cmult[44]) = (0,0);
		(Amult[30] => Cmult[44]) = (0,0);
		(Amult[31] => Cmult[44]) = (0,0);
		(Bmult[0]  => Cmult[44]) = (0,0);
		(Bmult[1]  => Cmult[44]) = (0,0);
		(Bmult[2]  => Cmult[44]) = (0,0);
		(Bmult[3]  => Cmult[44]) = (0,0);
		(Bmult[4]  => Cmult[44]) = (0,0);
		(Bmult[5]  => Cmult[44]) = (0,0);
		(Bmult[6]  => Cmult[44]) = (0,0);
		(Bmult[7]  => Cmult[44]) = (0,0);
		(Bmult[8]  => Cmult[44]) = (0,0);
		(Bmult[9]  => Cmult[44]) = (0,0);
		(Bmult[10] => Cmult[44]) = (0,0);
		(Bmult[11] => Cmult[44]) = (0,0);
		(Bmult[12] => Cmult[44]) = (0,0);
		(Bmult[13] => Cmult[44]) = (0,0);
		(Bmult[14] => Cmult[44]) = (0,0);
		(Bmult[15] => Cmult[44]) = (0,0);
		(Bmult[16] => Cmult[44]) = (0,0);
		(Bmult[17] => Cmult[44]) = (0,0);
		(Bmult[18] => Cmult[44]) = (0,0);
		(Bmult[19] => Cmult[44]) = (0,0);
		(Bmult[20] => Cmult[44]) = (0,0);
		(Bmult[21] => Cmult[44]) = (0,0);
		(Bmult[22] => Cmult[44]) = (0,0);
		(Bmult[23] => Cmult[44]) = (0,0);
		(Bmult[24] => Cmult[44]) = (0,0);
		(Bmult[25] => Cmult[44]) = (0,0);
		(Bmult[26] => Cmult[44]) = (0,0);
		(Bmult[27] => Cmult[44]) = (0,0);
		(Bmult[28] => Cmult[44]) = (0,0);
		(Bmult[29] => Cmult[44]) = (0,0);
		(Bmult[30] => Cmult[44]) = (0,0);
		(Bmult[31] => Cmult[44]) = (0,0);		
		(Valid_mult[0] => Cmult[44]) = (0,0);
		(Valid_mult[1] => Cmult[44]) = (0,0);
		(sel_mul_32x32 => Cmult[44]) = (0,0);
		(Amult[0]  => Cmult[45]) = (0,0);
		(Amult[1]  => Cmult[45]) = (0,0);
		(Amult[2]  => Cmult[45]) = (0,0);
		(Amult[3]  => Cmult[45]) = (0,0);
		(Amult[4]  => Cmult[45]) = (0,0);
		(Amult[5]  => Cmult[45]) = (0,0);
		(Amult[6]  => Cmult[45]) = (0,0);
		(Amult[7]  => Cmult[45]) = (0,0);
		(Amult[8]  => Cmult[45]) = (0,0);
		(Amult[9]  => Cmult[45]) = (0,0);
		(Amult[10] => Cmult[45]) = (0,0);
		(Amult[11] => Cmult[45]) = (0,0);
		(Amult[12] => Cmult[45]) = (0,0);
		(Amult[13] => Cmult[45]) = (0,0);
		(Amult[14] => Cmult[45]) = (0,0);
		(Amult[15] => Cmult[45]) = (0,0);
		(Amult[16] => Cmult[45]) = (0,0);
		(Amult[17] => Cmult[45]) = (0,0);
		(Amult[18] => Cmult[45]) = (0,0);
		(Amult[19] => Cmult[45]) = (0,0);
		(Amult[20] => Cmult[45]) = (0,0);
		(Amult[21] => Cmult[45]) = (0,0);
		(Amult[22] => Cmult[45]) = (0,0);
		(Amult[23] => Cmult[45]) = (0,0);
		(Amult[24] => Cmult[45]) = (0,0);
		(Amult[25] => Cmult[45]) = (0,0);
		(Amult[26] => Cmult[45]) = (0,0);
		(Amult[27] => Cmult[45]) = (0,0);
		(Amult[28] => Cmult[45]) = (0,0);
		(Amult[29] => Cmult[45]) = (0,0);
		(Amult[30] => Cmult[45]) = (0,0);
		(Amult[31] => Cmult[45]) = (0,0);
		(Bmult[0]  => Cmult[45]) = (0,0);
		(Bmult[1]  => Cmult[45]) = (0,0);
		(Bmult[2]  => Cmult[45]) = (0,0);
		(Bmult[3]  => Cmult[45]) = (0,0);
		(Bmult[4]  => Cmult[45]) = (0,0);
		(Bmult[5]  => Cmult[45]) = (0,0);
		(Bmult[6]  => Cmult[45]) = (0,0);
		(Bmult[7]  => Cmult[45]) = (0,0);
		(Bmult[8]  => Cmult[45]) = (0,0);
		(Bmult[9]  => Cmult[45]) = (0,0);
		(Bmult[10] => Cmult[45]) = (0,0);
		(Bmult[11] => Cmult[45]) = (0,0);
		(Bmult[12] => Cmult[45]) = (0,0);
		(Bmult[13] => Cmult[45]) = (0,0);
		(Bmult[14] => Cmult[45]) = (0,0);
		(Bmult[15] => Cmult[45]) = (0,0);
		(Bmult[16] => Cmult[45]) = (0,0);
		(Bmult[17] => Cmult[45]) = (0,0);
		(Bmult[18] => Cmult[45]) = (0,0);
		(Bmult[19] => Cmult[45]) = (0,0);
		(Bmult[20] => Cmult[45]) = (0,0);
		(Bmult[21] => Cmult[45]) = (0,0);
		(Bmult[22] => Cmult[45]) = (0,0);
		(Bmult[23] => Cmult[45]) = (0,0);
		(Bmult[24] => Cmult[45]) = (0,0);
		(Bmult[25] => Cmult[45]) = (0,0);
		(Bmult[26] => Cmult[45]) = (0,0);
		(Bmult[27] => Cmult[45]) = (0,0);
		(Bmult[28] => Cmult[45]) = (0,0);
		(Bmult[29] => Cmult[45]) = (0,0);
		(Bmult[30] => Cmult[45]) = (0,0);
		(Bmult[31] => Cmult[45]) = (0,0);		
		(Valid_mult[0] => Cmult[45]) = (0,0);
		(Valid_mult[1] => Cmult[45]) = (0,0);
		(sel_mul_32x32 => Cmult[45]) = (0,0);
		(Amult[0]  => Cmult[46]) = (0,0);
		(Amult[1]  => Cmult[46]) = (0,0);
		(Amult[2]  => Cmult[46]) = (0,0);
		(Amult[3]  => Cmult[46]) = (0,0);
		(Amult[4]  => Cmult[46]) = (0,0);
		(Amult[5]  => Cmult[46]) = (0,0);
		(Amult[6]  => Cmult[46]) = (0,0);
		(Amult[7]  => Cmult[46]) = (0,0);
		(Amult[8]  => Cmult[46]) = (0,0);
		(Amult[9]  => Cmult[46]) = (0,0);
		(Amult[10] => Cmult[46]) = (0,0);
		(Amult[11] => Cmult[46]) = (0,0);
		(Amult[12] => Cmult[46]) = (0,0);
		(Amult[13] => Cmult[46]) = (0,0);
		(Amult[14] => Cmult[46]) = (0,0);
		(Amult[15] => Cmult[46]) = (0,0);
		(Amult[16] => Cmult[46]) = (0,0);
		(Amult[17] => Cmult[46]) = (0,0);
		(Amult[18] => Cmult[46]) = (0,0);
		(Amult[19] => Cmult[46]) = (0,0);
		(Amult[20] => Cmult[46]) = (0,0);
		(Amult[21] => Cmult[46]) = (0,0);
		(Amult[22] => Cmult[46]) = (0,0);
		(Amult[23] => Cmult[46]) = (0,0);
		(Amult[24] => Cmult[46]) = (0,0);
		(Amult[25] => Cmult[46]) = (0,0);
		(Amult[26] => Cmult[46]) = (0,0);
		(Amult[27] => Cmult[46]) = (0,0);
		(Amult[28] => Cmult[46]) = (0,0);
		(Amult[29] => Cmult[46]) = (0,0);
		(Amult[30] => Cmult[46]) = (0,0);
		(Amult[31] => Cmult[46]) = (0,0);
		(Bmult[0]  => Cmult[46]) = (0,0);
		(Bmult[1]  => Cmult[46]) = (0,0);
		(Bmult[2]  => Cmult[46]) = (0,0);
		(Bmult[3]  => Cmult[46]) = (0,0);
		(Bmult[4]  => Cmult[46]) = (0,0);
		(Bmult[5]  => Cmult[46]) = (0,0);
		(Bmult[6]  => Cmult[46]) = (0,0);
		(Bmult[7]  => Cmult[46]) = (0,0);
		(Bmult[8]  => Cmult[46]) = (0,0);
		(Bmult[9]  => Cmult[46]) = (0,0);
		(Bmult[10] => Cmult[46]) = (0,0);
		(Bmult[11] => Cmult[46]) = (0,0);
		(Bmult[12] => Cmult[46]) = (0,0);
		(Bmult[13] => Cmult[46]) = (0,0);
		(Bmult[14] => Cmult[46]) = (0,0);
		(Bmult[15] => Cmult[46]) = (0,0);
		(Bmult[16] => Cmult[46]) = (0,0);
		(Bmult[17] => Cmult[46]) = (0,0);
		(Bmult[18] => Cmult[46]) = (0,0);
		(Bmult[19] => Cmult[46]) = (0,0);
		(Bmult[20] => Cmult[46]) = (0,0);
		(Bmult[21] => Cmult[46]) = (0,0);
		(Bmult[22] => Cmult[46]) = (0,0);
		(Bmult[23] => Cmult[46]) = (0,0);
		(Bmult[24] => Cmult[46]) = (0,0);
		(Bmult[25] => Cmult[46]) = (0,0);
		(Bmult[26] => Cmult[46]) = (0,0);
		(Bmult[27] => Cmult[46]) = (0,0);
		(Bmult[28] => Cmult[46]) = (0,0);
		(Bmult[29] => Cmult[46]) = (0,0);
		(Bmult[30] => Cmult[46]) = (0,0);
		(Bmult[31] => Cmult[46]) = (0,0);		
		(Valid_mult[0] => Cmult[46]) = (0,0);
		(Valid_mult[1] => Cmult[46]) = (0,0);
		(sel_mul_32x32 => Cmult[46]) = (0,0);
		(Amult[0]  => Cmult[47]) = (0,0);
		(Amult[1]  => Cmult[47]) = (0,0);
		(Amult[2]  => Cmult[47]) = (0,0);
		(Amult[3]  => Cmult[47]) = (0,0);
		(Amult[4]  => Cmult[47]) = (0,0);
		(Amult[5]  => Cmult[47]) = (0,0);
		(Amult[6]  => Cmult[47]) = (0,0);
		(Amult[7]  => Cmult[47]) = (0,0);
		(Amult[8]  => Cmult[47]) = (0,0);
		(Amult[9]  => Cmult[47]) = (0,0);
		(Amult[10] => Cmult[47]) = (0,0);
		(Amult[11] => Cmult[47]) = (0,0);
		(Amult[12] => Cmult[47]) = (0,0);
		(Amult[13] => Cmult[47]) = (0,0);
		(Amult[14] => Cmult[47]) = (0,0);
		(Amult[15] => Cmult[47]) = (0,0);
		(Amult[16] => Cmult[47]) = (0,0);
		(Amult[17] => Cmult[47]) = (0,0);
		(Amult[18] => Cmult[47]) = (0,0);
		(Amult[19] => Cmult[47]) = (0,0);
		(Amult[20] => Cmult[47]) = (0,0);
		(Amult[21] => Cmult[47]) = (0,0);
		(Amult[22] => Cmult[47]) = (0,0);
		(Amult[23] => Cmult[47]) = (0,0);
		(Amult[24] => Cmult[47]) = (0,0);
		(Amult[25] => Cmult[47]) = (0,0);
		(Amult[26] => Cmult[47]) = (0,0);
		(Amult[27] => Cmult[47]) = (0,0);
		(Amult[28] => Cmult[47]) = (0,0);
		(Amult[29] => Cmult[47]) = (0,0);
		(Amult[30] => Cmult[47]) = (0,0);
		(Amult[31] => Cmult[47]) = (0,0);
		(Bmult[0]  => Cmult[47]) = (0,0);
		(Bmult[1]  => Cmult[47]) = (0,0);
		(Bmult[2]  => Cmult[47]) = (0,0);
		(Bmult[3]  => Cmult[47]) = (0,0);
		(Bmult[4]  => Cmult[47]) = (0,0);
		(Bmult[5]  => Cmult[47]) = (0,0);
		(Bmult[6]  => Cmult[47]) = (0,0);
		(Bmult[7]  => Cmult[47]) = (0,0);
		(Bmult[8]  => Cmult[47]) = (0,0);
		(Bmult[9]  => Cmult[47]) = (0,0);
		(Bmult[10] => Cmult[47]) = (0,0);
		(Bmult[11] => Cmult[47]) = (0,0);
		(Bmult[12] => Cmult[47]) = (0,0);
		(Bmult[13] => Cmult[47]) = (0,0);
		(Bmult[14] => Cmult[47]) = (0,0);
		(Bmult[15] => Cmult[47]) = (0,0);
		(Bmult[16] => Cmult[47]) = (0,0);
		(Bmult[17] => Cmult[47]) = (0,0);
		(Bmult[18] => Cmult[47]) = (0,0);
		(Bmult[19] => Cmult[47]) = (0,0);
		(Bmult[20] => Cmult[47]) = (0,0);
		(Bmult[21] => Cmult[47]) = (0,0);
		(Bmult[22] => Cmult[47]) = (0,0);
		(Bmult[23] => Cmult[47]) = (0,0);
		(Bmult[24] => Cmult[47]) = (0,0);
		(Bmult[25] => Cmult[47]) = (0,0);
		(Bmult[26] => Cmult[47]) = (0,0);
		(Bmult[27] => Cmult[47]) = (0,0);
		(Bmult[28] => Cmult[47]) = (0,0);
		(Bmult[29] => Cmult[47]) = (0,0);
		(Bmult[30] => Cmult[47]) = (0,0);
		(Bmult[31] => Cmult[47]) = (0,0);		
		(Valid_mult[0] => Cmult[47]) = (0,0);
		(Valid_mult[1] => Cmult[47]) = (0,0);
		(sel_mul_32x32 => Cmult[47]) = (0,0);
		(Amult[0]  => Cmult[48]) = (0,0);
		(Amult[1]  => Cmult[48]) = (0,0);
		(Amult[2]  => Cmult[48]) = (0,0);
		(Amult[3]  => Cmult[48]) = (0,0);
		(Amult[4]  => Cmult[48]) = (0,0);
		(Amult[5]  => Cmult[48]) = (0,0);
		(Amult[6]  => Cmult[48]) = (0,0);
		(Amult[7]  => Cmult[48]) = (0,0);
		(Amult[8]  => Cmult[48]) = (0,0);
		(Amult[9]  => Cmult[48]) = (0,0);
		(Amult[10] => Cmult[48]) = (0,0);
		(Amult[11] => Cmult[48]) = (0,0);
		(Amult[12] => Cmult[48]) = (0,0);
		(Amult[13] => Cmult[48]) = (0,0);
		(Amult[14] => Cmult[48]) = (0,0);
		(Amult[15] => Cmult[48]) = (0,0);
		(Amult[16] => Cmult[48]) = (0,0);
		(Amult[17] => Cmult[48]) = (0,0);
		(Amult[18] => Cmult[48]) = (0,0);
		(Amult[19] => Cmult[48]) = (0,0);
		(Amult[20] => Cmult[48]) = (0,0);
		(Amult[21] => Cmult[48]) = (0,0);
		(Amult[22] => Cmult[48]) = (0,0);
		(Amult[23] => Cmult[48]) = (0,0);
		(Amult[24] => Cmult[48]) = (0,0);
		(Amult[25] => Cmult[48]) = (0,0);
		(Amult[26] => Cmult[48]) = (0,0);
		(Amult[27] => Cmult[48]) = (0,0);
		(Amult[28] => Cmult[48]) = (0,0);
		(Amult[29] => Cmult[48]) = (0,0);
		(Amult[30] => Cmult[48]) = (0,0);
		(Amult[31] => Cmult[48]) = (0,0);
		(Bmult[0]  => Cmult[48]) = (0,0);
		(Bmult[1]  => Cmult[48]) = (0,0);
		(Bmult[2]  => Cmult[48]) = (0,0);
		(Bmult[3]  => Cmult[48]) = (0,0);
		(Bmult[4]  => Cmult[48]) = (0,0);
		(Bmult[5]  => Cmult[48]) = (0,0);
		(Bmult[6]  => Cmult[48]) = (0,0);
		(Bmult[7]  => Cmult[48]) = (0,0);
		(Bmult[8]  => Cmult[48]) = (0,0);
		(Bmult[9]  => Cmult[48]) = (0,0);
		(Bmult[10] => Cmult[48]) = (0,0);
		(Bmult[11] => Cmult[48]) = (0,0);
		(Bmult[12] => Cmult[48]) = (0,0);
		(Bmult[13] => Cmult[48]) = (0,0);
		(Bmult[14] => Cmult[48]) = (0,0);
		(Bmult[15] => Cmult[48]) = (0,0);
		(Bmult[16] => Cmult[48]) = (0,0);
		(Bmult[17] => Cmult[48]) = (0,0);
		(Bmult[18] => Cmult[48]) = (0,0);
		(Bmult[19] => Cmult[48]) = (0,0);
		(Bmult[20] => Cmult[48]) = (0,0);
		(Bmult[21] => Cmult[48]) = (0,0);
		(Bmult[22] => Cmult[48]) = (0,0);
		(Bmult[23] => Cmult[48]) = (0,0);
		(Bmult[24] => Cmult[48]) = (0,0);
		(Bmult[25] => Cmult[48]) = (0,0);
		(Bmult[26] => Cmult[48]) = (0,0);
		(Bmult[27] => Cmult[48]) = (0,0);
		(Bmult[28] => Cmult[48]) = (0,0);
		(Bmult[29] => Cmult[48]) = (0,0);
		(Bmult[30] => Cmult[48]) = (0,0);
		(Bmult[31] => Cmult[48]) = (0,0);		
		(Valid_mult[0] => Cmult[48]) = (0,0);
		(Valid_mult[1] => Cmult[48]) = (0,0);
		(sel_mul_32x32 => Cmult[48]) = (0,0);	
		(Amult[0]  => Cmult[49]) = (0,0);
		(Amult[1]  => Cmult[49]) = (0,0);
		(Amult[2]  => Cmult[49]) = (0,0);
		(Amult[3]  => Cmult[49]) = (0,0);
		(Amult[4]  => Cmult[49]) = (0,0);
		(Amult[5]  => Cmult[49]) = (0,0);
		(Amult[6]  => Cmult[49]) = (0,0);
		(Amult[7]  => Cmult[49]) = (0,0);
		(Amult[8]  => Cmult[49]) = (0,0);
		(Amult[9]  => Cmult[49]) = (0,0);
		(Amult[10] => Cmult[49]) = (0,0);
		(Amult[11] => Cmult[49]) = (0,0);
		(Amult[12] => Cmult[49]) = (0,0);
		(Amult[13] => Cmult[49]) = (0,0);
		(Amult[14] => Cmult[49]) = (0,0);
		(Amult[15] => Cmult[49]) = (0,0);
		(Amult[16] => Cmult[49]) = (0,0);
		(Amult[17] => Cmult[49]) = (0,0);
		(Amult[18] => Cmult[49]) = (0,0);
		(Amult[19] => Cmult[49]) = (0,0);
		(Amult[20] => Cmult[49]) = (0,0);
		(Amult[21] => Cmult[49]) = (0,0);
		(Amult[22] => Cmult[49]) = (0,0);
		(Amult[23] => Cmult[49]) = (0,0);
		(Amult[24] => Cmult[49]) = (0,0);
		(Amult[25] => Cmult[49]) = (0,0);
		(Amult[26] => Cmult[49]) = (0,0);
		(Amult[27] => Cmult[49]) = (0,0);
		(Amult[28] => Cmult[49]) = (0,0);
		(Amult[29] => Cmult[49]) = (0,0);
		(Amult[30] => Cmult[49]) = (0,0);
		(Amult[31] => Cmult[49]) = (0,0);
		(Bmult[0]  => Cmult[49]) = (0,0);
		(Bmult[1]  => Cmult[49]) = (0,0);
		(Bmult[2]  => Cmult[49]) = (0,0);
		(Bmult[3]  => Cmult[49]) = (0,0);
		(Bmult[4]  => Cmult[49]) = (0,0);
		(Bmult[5]  => Cmult[49]) = (0,0);
		(Bmult[6]  => Cmult[49]) = (0,0);
		(Bmult[7]  => Cmult[49]) = (0,0);
		(Bmult[8]  => Cmult[49]) = (0,0);
		(Bmult[9]  => Cmult[49]) = (0,0);
		(Bmult[10] => Cmult[49]) = (0,0);
		(Bmult[11] => Cmult[49]) = (0,0);
		(Bmult[12] => Cmult[49]) = (0,0);
		(Bmult[13] => Cmult[49]) = (0,0);
		(Bmult[14] => Cmult[49]) = (0,0);
		(Bmult[15] => Cmult[49]) = (0,0);
		(Bmult[16] => Cmult[49]) = (0,0);
		(Bmult[17] => Cmult[49]) = (0,0);
		(Bmult[18] => Cmult[49]) = (0,0);
		(Bmult[19] => Cmult[49]) = (0,0);
		(Bmult[20] => Cmult[49]) = (0,0);
		(Bmult[21] => Cmult[49]) = (0,0);
		(Bmult[22] => Cmult[49]) = (0,0);
		(Bmult[23] => Cmult[49]) = (0,0);
		(Bmult[24] => Cmult[49]) = (0,0);
		(Bmult[25] => Cmult[49]) = (0,0);
		(Bmult[26] => Cmult[49]) = (0,0);
		(Bmult[27] => Cmult[49]) = (0,0);
		(Bmult[28] => Cmult[49]) = (0,0);
		(Bmult[29] => Cmult[49]) = (0,0);
		(Bmult[30] => Cmult[49]) = (0,0);
		(Bmult[31] => Cmult[49]) = (0,0);		
		(Valid_mult[0] => Cmult[49]) = (0,0);
		(Valid_mult[1] => Cmult[49]) = (0,0);
		(sel_mul_32x32 => Cmult[49]) = (0,0);
		(Amult[0]  => Cmult[50]) = (0,0);
		(Amult[1]  => Cmult[50]) = (0,0);
		(Amult[2]  => Cmult[50]) = (0,0);
		(Amult[3]  => Cmult[50]) = (0,0);
		(Amult[4]  => Cmult[50]) = (0,0);
		(Amult[5]  => Cmult[50]) = (0,0);
		(Amult[6]  => Cmult[50]) = (0,0);
		(Amult[7]  => Cmult[50]) = (0,0);
		(Amult[8]  => Cmult[50]) = (0,0);
		(Amult[9]  => Cmult[50]) = (0,0);
		(Amult[10] => Cmult[50]) = (0,0);
		(Amult[11] => Cmult[50]) = (0,0);
		(Amult[12] => Cmult[50]) = (0,0);
		(Amult[13] => Cmult[50]) = (0,0);
		(Amult[14] => Cmult[50]) = (0,0);
		(Amult[15] => Cmult[50]) = (0,0);
		(Amult[16] => Cmult[50]) = (0,0);
		(Amult[17] => Cmult[50]) = (0,0);
		(Amult[18] => Cmult[50]) = (0,0);
		(Amult[19] => Cmult[50]) = (0,0);
		(Amult[20] => Cmult[50]) = (0,0);
		(Amult[21] => Cmult[50]) = (0,0);
		(Amult[22] => Cmult[50]) = (0,0);
		(Amult[23] => Cmult[50]) = (0,0);
		(Amult[24] => Cmult[50]) = (0,0);
		(Amult[25] => Cmult[50]) = (0,0);
		(Amult[26] => Cmult[50]) = (0,0);
		(Amult[27] => Cmult[50]) = (0,0);
		(Amult[28] => Cmult[50]) = (0,0);
		(Amult[29] => Cmult[50]) = (0,0);
		(Amult[30] => Cmult[50]) = (0,0);
		(Amult[31] => Cmult[50]) = (0,0);
		(Bmult[0]  => Cmult[50]) = (0,0);
		(Bmult[1]  => Cmult[50]) = (0,0);
		(Bmult[2]  => Cmult[50]) = (0,0);
		(Bmult[3]  => Cmult[50]) = (0,0);
		(Bmult[4]  => Cmult[50]) = (0,0);
		(Bmult[5]  => Cmult[50]) = (0,0);
		(Bmult[6]  => Cmult[50]) = (0,0);
		(Bmult[7]  => Cmult[50]) = (0,0);
		(Bmult[8]  => Cmult[50]) = (0,0);
		(Bmult[9]  => Cmult[50]) = (0,0);
		(Bmult[10] => Cmult[50]) = (0,0);
		(Bmult[11] => Cmult[50]) = (0,0);
		(Bmult[12] => Cmult[50]) = (0,0);
		(Bmult[13] => Cmult[50]) = (0,0);
		(Bmult[14] => Cmult[50]) = (0,0);
		(Bmult[15] => Cmult[50]) = (0,0);
		(Bmult[16] => Cmult[50]) = (0,0);
		(Bmult[17] => Cmult[50]) = (0,0);
		(Bmult[18] => Cmult[50]) = (0,0);
		(Bmult[19] => Cmult[50]) = (0,0);
		(Bmult[20] => Cmult[50]) = (0,0);
		(Bmult[21] => Cmult[50]) = (0,0);
		(Bmult[22] => Cmult[50]) = (0,0);
		(Bmult[23] => Cmult[50]) = (0,0);
		(Bmult[24] => Cmult[50]) = (0,0);
		(Bmult[25] => Cmult[50]) = (0,0);
		(Bmult[26] => Cmult[50]) = (0,0);
		(Bmult[27] => Cmult[50]) = (0,0);
		(Bmult[28] => Cmult[50]) = (0,0);
		(Bmult[29] => Cmult[50]) = (0,0);
		(Bmult[30] => Cmult[50]) = (0,0);
		(Bmult[31] => Cmult[50]) = (0,0);		
		(Valid_mult[0] => Cmult[50]) = (0,0);
		(Valid_mult[1] => Cmult[50]) = (0,0);
		(sel_mul_32x32 => Cmult[50]) = (0,0);
		(Amult[0]  => Cmult[51]) = (0,0);
		(Amult[1]  => Cmult[51]) = (0,0);
		(Amult[2]  => Cmult[51]) = (0,0);
		(Amult[3]  => Cmult[51]) = (0,0);
		(Amult[4]  => Cmult[51]) = (0,0);
		(Amult[5]  => Cmult[51]) = (0,0);
		(Amult[6]  => Cmult[51]) = (0,0);
		(Amult[7]  => Cmult[51]) = (0,0);
		(Amult[8]  => Cmult[51]) = (0,0);
		(Amult[9]  => Cmult[51]) = (0,0);
		(Amult[10] => Cmult[51]) = (0,0);
		(Amult[11] => Cmult[51]) = (0,0);
		(Amult[12] => Cmult[51]) = (0,0);
		(Amult[13] => Cmult[51]) = (0,0);
		(Amult[14] => Cmult[51]) = (0,0);
		(Amult[15] => Cmult[51]) = (0,0);
		(Amult[16] => Cmult[51]) = (0,0);
		(Amult[17] => Cmult[51]) = (0,0);
		(Amult[18] => Cmult[51]) = (0,0);
		(Amult[19] => Cmult[51]) = (0,0);
		(Amult[20] => Cmult[51]) = (0,0);
		(Amult[21] => Cmult[51]) = (0,0);
		(Amult[22] => Cmult[51]) = (0,0);
		(Amult[23] => Cmult[51]) = (0,0);
		(Amult[24] => Cmult[51]) = (0,0);
		(Amult[25] => Cmult[51]) = (0,0);
		(Amult[26] => Cmult[51]) = (0,0);
		(Amult[27] => Cmult[51]) = (0,0);
		(Amult[28] => Cmult[51]) = (0,0);
		(Amult[29] => Cmult[51]) = (0,0);
		(Amult[30] => Cmult[51]) = (0,0);
		(Amult[31] => Cmult[51]) = (0,0);
		(Bmult[0]  => Cmult[51]) = (0,0);
		(Bmult[1]  => Cmult[51]) = (0,0);
		(Bmult[2]  => Cmult[51]) = (0,0);
		(Bmult[3]  => Cmult[51]) = (0,0);
		(Bmult[4]  => Cmult[51]) = (0,0);
		(Bmult[5]  => Cmult[51]) = (0,0);
		(Bmult[6]  => Cmult[51]) = (0,0);
		(Bmult[7]  => Cmult[51]) = (0,0);
		(Bmult[8]  => Cmult[51]) = (0,0);
		(Bmult[9]  => Cmult[51]) = (0,0);
		(Bmult[10] => Cmult[51]) = (0,0);
		(Bmult[11] => Cmult[51]) = (0,0);
		(Bmult[12] => Cmult[51]) = (0,0);
		(Bmult[13] => Cmult[51]) = (0,0);
		(Bmult[14] => Cmult[51]) = (0,0);
		(Bmult[15] => Cmult[51]) = (0,0);
		(Bmult[16] => Cmult[51]) = (0,0);
		(Bmult[17] => Cmult[51]) = (0,0);
		(Bmult[18] => Cmult[51]) = (0,0);
		(Bmult[19] => Cmult[51]) = (0,0);
		(Bmult[20] => Cmult[51]) = (0,0);
		(Bmult[21] => Cmult[51]) = (0,0);
		(Bmult[22] => Cmult[51]) = (0,0);
		(Bmult[23] => Cmult[51]) = (0,0);
		(Bmult[24] => Cmult[51]) = (0,0);
		(Bmult[25] => Cmult[51]) = (0,0);
		(Bmult[26] => Cmult[51]) = (0,0);
		(Bmult[27] => Cmult[51]) = (0,0);
		(Bmult[28] => Cmult[51]) = (0,0);
		(Bmult[29] => Cmult[51]) = (0,0);
		(Bmult[30] => Cmult[51]) = (0,0);
		(Bmult[31] => Cmult[51]) = (0,0);		
		(Valid_mult[0] => Cmult[51]) = (0,0);
		(Valid_mult[1] => Cmult[51]) = (0,0);
		(sel_mul_32x32 => Cmult[51]) = (0,0);
		(Amult[0]  => Cmult[52]) = (0,0);
		(Amult[1]  => Cmult[52]) = (0,0);
		(Amult[2]  => Cmult[52]) = (0,0);
		(Amult[3]  => Cmult[52]) = (0,0);
		(Amult[4]  => Cmult[52]) = (0,0);
		(Amult[5]  => Cmult[52]) = (0,0);
		(Amult[6]  => Cmult[52]) = (0,0);
		(Amult[7]  => Cmult[52]) = (0,0);
		(Amult[8]  => Cmult[52]) = (0,0);
		(Amult[9]  => Cmult[52]) = (0,0);
		(Amult[10] => Cmult[52]) = (0,0);
		(Amult[11] => Cmult[52]) = (0,0);
		(Amult[12] => Cmult[52]) = (0,0);
		(Amult[13] => Cmult[52]) = (0,0);
		(Amult[14] => Cmult[52]) = (0,0);
		(Amult[15] => Cmult[52]) = (0,0);
		(Amult[16] => Cmult[52]) = (0,0);
		(Amult[17] => Cmult[52]) = (0,0);
		(Amult[18] => Cmult[52]) = (0,0);
		(Amult[19] => Cmult[52]) = (0,0);
		(Amult[20] => Cmult[52]) = (0,0);
		(Amult[21] => Cmult[52]) = (0,0);
		(Amult[22] => Cmult[52]) = (0,0);
		(Amult[23] => Cmult[52]) = (0,0);
		(Amult[24] => Cmult[52]) = (0,0);
		(Amult[25] => Cmult[52]) = (0,0);
		(Amult[26] => Cmult[52]) = (0,0);
		(Amult[27] => Cmult[52]) = (0,0);
		(Amult[28] => Cmult[52]) = (0,0);
		(Amult[29] => Cmult[52]) = (0,0);
		(Amult[30] => Cmult[52]) = (0,0);
		(Amult[31] => Cmult[52]) = (0,0);
		(Bmult[0]  => Cmult[52]) = (0,0);
		(Bmult[1]  => Cmult[52]) = (0,0);
		(Bmult[2]  => Cmult[52]) = (0,0);
		(Bmult[3]  => Cmult[52]) = (0,0);
		(Bmult[4]  => Cmult[52]) = (0,0);
		(Bmult[5]  => Cmult[52]) = (0,0);
		(Bmult[6]  => Cmult[52]) = (0,0);
		(Bmult[7]  => Cmult[52]) = (0,0);
		(Bmult[8]  => Cmult[52]) = (0,0);
		(Bmult[9]  => Cmult[52]) = (0,0);
		(Bmult[10] => Cmult[52]) = (0,0);
		(Bmult[11] => Cmult[52]) = (0,0);
		(Bmult[12] => Cmult[52]) = (0,0);
		(Bmult[13] => Cmult[52]) = (0,0);
		(Bmult[14] => Cmult[52]) = (0,0);
		(Bmult[15] => Cmult[52]) = (0,0);
		(Bmult[16] => Cmult[52]) = (0,0);
		(Bmult[17] => Cmult[52]) = (0,0);
		(Bmult[18] => Cmult[52]) = (0,0);
		(Bmult[19] => Cmult[52]) = (0,0);
		(Bmult[20] => Cmult[52]) = (0,0);
		(Bmult[21] => Cmult[52]) = (0,0);
		(Bmult[22] => Cmult[52]) = (0,0);
		(Bmult[23] => Cmult[52]) = (0,0);
		(Bmult[24] => Cmult[52]) = (0,0);
		(Bmult[25] => Cmult[52]) = (0,0);
		(Bmult[26] => Cmult[52]) = (0,0);
		(Bmult[27] => Cmult[52]) = (0,0);
		(Bmult[28] => Cmult[52]) = (0,0);
		(Bmult[29] => Cmult[52]) = (0,0);
		(Bmult[30] => Cmult[52]) = (0,0);
		(Bmult[31] => Cmult[52]) = (0,0);		
		(Valid_mult[0] => Cmult[52]) = (0,0);
		(Valid_mult[1] => Cmult[52]) = (0,0);
		(sel_mul_32x32 => Cmult[52]) = (0,0);
		(Amult[0]  => Cmult[53]) = (0,0);
		(Amult[1]  => Cmult[53]) = (0,0);
		(Amult[2]  => Cmult[53]) = (0,0);
		(Amult[3]  => Cmult[53]) = (0,0);
		(Amult[4]  => Cmult[53]) = (0,0);
		(Amult[5]  => Cmult[53]) = (0,0);
		(Amult[6]  => Cmult[53]) = (0,0);
		(Amult[7]  => Cmult[53]) = (0,0);
		(Amult[8]  => Cmult[53]) = (0,0);
		(Amult[9]  => Cmult[53]) = (0,0);
		(Amult[10] => Cmult[53]) = (0,0);
		(Amult[11] => Cmult[53]) = (0,0);
		(Amult[12] => Cmult[53]) = (0,0);
		(Amult[13] => Cmult[53]) = (0,0);
		(Amult[14] => Cmult[53]) = (0,0);
		(Amult[15] => Cmult[53]) = (0,0);
		(Amult[16] => Cmult[53]) = (0,0);
		(Amult[17] => Cmult[53]) = (0,0);
		(Amult[18] => Cmult[53]) = (0,0);
		(Amult[19] => Cmult[53]) = (0,0);
		(Amult[20] => Cmult[53]) = (0,0);
		(Amult[21] => Cmult[53]) = (0,0);
		(Amult[22] => Cmult[53]) = (0,0);
		(Amult[23] => Cmult[53]) = (0,0);
		(Amult[24] => Cmult[53]) = (0,0);
		(Amult[25] => Cmult[53]) = (0,0);
		(Amult[26] => Cmult[53]) = (0,0);
		(Amult[27] => Cmult[53]) = (0,0);
		(Amult[28] => Cmult[53]) = (0,0);
		(Amult[29] => Cmult[53]) = (0,0);
		(Amult[30] => Cmult[53]) = (0,0);
		(Amult[31] => Cmult[53]) = (0,0);
		(Bmult[0]  => Cmult[53]) = (0,0);
		(Bmult[1]  => Cmult[53]) = (0,0);
		(Bmult[2]  => Cmult[53]) = (0,0);
		(Bmult[3]  => Cmult[53]) = (0,0);
		(Bmult[4]  => Cmult[53]) = (0,0);
		(Bmult[5]  => Cmult[53]) = (0,0);
		(Bmult[6]  => Cmult[53]) = (0,0);
		(Bmult[7]  => Cmult[53]) = (0,0);
		(Bmult[8]  => Cmult[53]) = (0,0);
		(Bmult[9]  => Cmult[53]) = (0,0);
		(Bmult[10] => Cmult[53]) = (0,0);
		(Bmult[11] => Cmult[53]) = (0,0);
		(Bmult[12] => Cmult[53]) = (0,0);
		(Bmult[13] => Cmult[53]) = (0,0);
		(Bmult[14] => Cmult[53]) = (0,0);
		(Bmult[15] => Cmult[53]) = (0,0);
		(Bmult[16] => Cmult[53]) = (0,0);
		(Bmult[17] => Cmult[53]) = (0,0);
		(Bmult[18] => Cmult[53]) = (0,0);
		(Bmult[19] => Cmult[53]) = (0,0);
		(Bmult[20] => Cmult[53]) = (0,0);
		(Bmult[21] => Cmult[53]) = (0,0);
		(Bmult[22] => Cmult[53]) = (0,0);
		(Bmult[23] => Cmult[53]) = (0,0);
		(Bmult[24] => Cmult[53]) = (0,0);
		(Bmult[25] => Cmult[53]) = (0,0);
		(Bmult[26] => Cmult[53]) = (0,0);
		(Bmult[27] => Cmult[53]) = (0,0);
		(Bmult[28] => Cmult[53]) = (0,0);
		(Bmult[29] => Cmult[53]) = (0,0);
		(Bmult[30] => Cmult[53]) = (0,0);
		(Bmult[31] => Cmult[53]) = (0,0);		
		(Valid_mult[0] => Cmult[53]) = (0,0);
		(Valid_mult[1] => Cmult[53]) = (0,0);
		(sel_mul_32x32 => Cmult[53]) = (0,0);
		(Amult[0]  => Cmult[54]) = (0,0);
		(Amult[1]  => Cmult[54]) = (0,0);
		(Amult[2]  => Cmult[54]) = (0,0);
		(Amult[3]  => Cmult[54]) = (0,0);
		(Amult[4]  => Cmult[54]) = (0,0);
		(Amult[5]  => Cmult[54]) = (0,0);
		(Amult[6]  => Cmult[54]) = (0,0);
		(Amult[7]  => Cmult[54]) = (0,0);
		(Amult[8]  => Cmult[54]) = (0,0);
		(Amult[9]  => Cmult[54]) = (0,0);
		(Amult[10] => Cmult[54]) = (0,0);
		(Amult[11] => Cmult[54]) = (0,0);
		(Amult[12] => Cmult[54]) = (0,0);
		(Amult[13] => Cmult[54]) = (0,0);
		(Amult[14] => Cmult[54]) = (0,0);
		(Amult[15] => Cmult[54]) = (0,0);
		(Amult[16] => Cmult[54]) = (0,0);
		(Amult[17] => Cmult[54]) = (0,0);
		(Amult[18] => Cmult[54]) = (0,0);
		(Amult[19] => Cmult[54]) = (0,0);
		(Amult[20] => Cmult[54]) = (0,0);
		(Amult[21] => Cmult[54]) = (0,0);
		(Amult[22] => Cmult[54]) = (0,0);
		(Amult[23] => Cmult[54]) = (0,0);
		(Amult[24] => Cmult[54]) = (0,0);
		(Amult[25] => Cmult[54]) = (0,0);
		(Amult[26] => Cmult[54]) = (0,0);
		(Amult[27] => Cmult[54]) = (0,0);
		(Amult[28] => Cmult[54]) = (0,0);
		(Amult[29] => Cmult[54]) = (0,0);
		(Amult[30] => Cmult[54]) = (0,0);
		(Amult[31] => Cmult[54]) = (0,0);
		(Bmult[0]  => Cmult[54]) = (0,0);
		(Bmult[1]  => Cmult[54]) = (0,0);
		(Bmult[2]  => Cmult[54]) = (0,0);
		(Bmult[3]  => Cmult[54]) = (0,0);
		(Bmult[4]  => Cmult[54]) = (0,0);
		(Bmult[5]  => Cmult[54]) = (0,0);
		(Bmult[6]  => Cmult[54]) = (0,0);
		(Bmult[7]  => Cmult[54]) = (0,0);
		(Bmult[8]  => Cmult[54]) = (0,0);
		(Bmult[9]  => Cmult[54]) = (0,0);
		(Bmult[10] => Cmult[54]) = (0,0);
		(Bmult[11] => Cmult[54]) = (0,0);
		(Bmult[12] => Cmult[54]) = (0,0);
		(Bmult[13] => Cmult[54]) = (0,0);
		(Bmult[14] => Cmult[54]) = (0,0);
		(Bmult[15] => Cmult[54]) = (0,0);
		(Bmult[16] => Cmult[54]) = (0,0);
		(Bmult[17] => Cmult[54]) = (0,0);
		(Bmult[18] => Cmult[54]) = (0,0);
		(Bmult[19] => Cmult[54]) = (0,0);
		(Bmult[20] => Cmult[54]) = (0,0);
		(Bmult[21] => Cmult[54]) = (0,0);
		(Bmult[22] => Cmult[54]) = (0,0);
		(Bmult[23] => Cmult[54]) = (0,0);
		(Bmult[24] => Cmult[54]) = (0,0);
		(Bmult[25] => Cmult[54]) = (0,0);
		(Bmult[26] => Cmult[54]) = (0,0);
		(Bmult[27] => Cmult[54]) = (0,0);
		(Bmult[28] => Cmult[54]) = (0,0);
		(Bmult[29] => Cmult[54]) = (0,0);
		(Bmult[30] => Cmult[54]) = (0,0);
		(Bmult[31] => Cmult[54]) = (0,0);		
		(Valid_mult[0] => Cmult[54]) = (0,0);
		(Valid_mult[1] => Cmult[54]) = (0,0);
		(sel_mul_32x32 => Cmult[54]) = (0,0);
		(Amult[0]  => Cmult[55]) = (0,0);
		(Amult[1]  => Cmult[55]) = (0,0);
		(Amult[2]  => Cmult[55]) = (0,0);
		(Amult[3]  => Cmult[55]) = (0,0);
		(Amult[4]  => Cmult[55]) = (0,0);
		(Amult[5]  => Cmult[55]) = (0,0);
		(Amult[6]  => Cmult[55]) = (0,0);
		(Amult[7]  => Cmult[55]) = (0,0);
		(Amult[8]  => Cmult[55]) = (0,0);
		(Amult[9]  => Cmult[55]) = (0,0);
		(Amult[10] => Cmult[55]) = (0,0);
		(Amult[11] => Cmult[55]) = (0,0);
		(Amult[12] => Cmult[55]) = (0,0);
		(Amult[13] => Cmult[55]) = (0,0);
		(Amult[14] => Cmult[55]) = (0,0);
		(Amult[15] => Cmult[55]) = (0,0);
		(Amult[16] => Cmult[55]) = (0,0);
		(Amult[17] => Cmult[55]) = (0,0);
		(Amult[18] => Cmult[55]) = (0,0);
		(Amult[19] => Cmult[55]) = (0,0);
		(Amult[20] => Cmult[55]) = (0,0);
		(Amult[21] => Cmult[55]) = (0,0);
		(Amult[22] => Cmult[55]) = (0,0);
		(Amult[23] => Cmult[55]) = (0,0);
		(Amult[24] => Cmult[55]) = (0,0);
		(Amult[25] => Cmult[55]) = (0,0);
		(Amult[26] => Cmult[55]) = (0,0);
		(Amult[27] => Cmult[55]) = (0,0);
		(Amult[28] => Cmult[55]) = (0,0);
		(Amult[29] => Cmult[55]) = (0,0);
		(Amult[30] => Cmult[55]) = (0,0);
		(Amult[31] => Cmult[55]) = (0,0);
		(Bmult[0]  => Cmult[55]) = (0,0);
		(Bmult[1]  => Cmult[55]) = (0,0);
		(Bmult[2]  => Cmult[55]) = (0,0);
		(Bmult[3]  => Cmult[55]) = (0,0);
		(Bmult[4]  => Cmult[55]) = (0,0);
		(Bmult[5]  => Cmult[55]) = (0,0);
		(Bmult[6]  => Cmult[55]) = (0,0);
		(Bmult[7]  => Cmult[55]) = (0,0);
		(Bmult[8]  => Cmult[55]) = (0,0);
		(Bmult[9]  => Cmult[55]) = (0,0);
		(Bmult[10] => Cmult[55]) = (0,0);
		(Bmult[11] => Cmult[55]) = (0,0);
		(Bmult[12] => Cmult[55]) = (0,0);
		(Bmult[13] => Cmult[55]) = (0,0);
		(Bmult[14] => Cmult[55]) = (0,0);
		(Bmult[15] => Cmult[55]) = (0,0);
		(Bmult[16] => Cmult[55]) = (0,0);
		(Bmult[17] => Cmult[55]) = (0,0);
		(Bmult[18] => Cmult[55]) = (0,0);
		(Bmult[19] => Cmult[55]) = (0,0);
		(Bmult[20] => Cmult[55]) = (0,0);
		(Bmult[21] => Cmult[55]) = (0,0);
		(Bmult[22] => Cmult[55]) = (0,0);
		(Bmult[23] => Cmult[55]) = (0,0);
		(Bmult[24] => Cmult[55]) = (0,0);
		(Bmult[25] => Cmult[55]) = (0,0);
		(Bmult[26] => Cmult[55]) = (0,0);
		(Bmult[27] => Cmult[55]) = (0,0);
		(Bmult[28] => Cmult[55]) = (0,0);
		(Bmult[29] => Cmult[55]) = (0,0);
		(Bmult[30] => Cmult[55]) = (0,0);
		(Bmult[31] => Cmult[55]) = (0,0);		
		(Valid_mult[0] => Cmult[55]) = (0,0);
		(Valid_mult[1] => Cmult[55]) = (0,0);
		(sel_mul_32x32 => Cmult[55]) = (0,0);
		(Amult[0]  => Cmult[56]) = (0,0);
		(Amult[1]  => Cmult[56]) = (0,0);
		(Amult[2]  => Cmult[56]) = (0,0);
		(Amult[3]  => Cmult[56]) = (0,0);
		(Amult[4]  => Cmult[56]) = (0,0);
		(Amult[5]  => Cmult[56]) = (0,0);
		(Amult[6]  => Cmult[56]) = (0,0);
		(Amult[7]  => Cmult[56]) = (0,0);
		(Amult[8]  => Cmult[56]) = (0,0);
		(Amult[9]  => Cmult[56]) = (0,0);
		(Amult[10] => Cmult[56]) = (0,0);
		(Amult[11] => Cmult[56]) = (0,0);
		(Amult[12] => Cmult[56]) = (0,0);
		(Amult[13] => Cmult[56]) = (0,0);
		(Amult[14] => Cmult[56]) = (0,0);
		(Amult[15] => Cmult[56]) = (0,0);
		(Amult[16] => Cmult[56]) = (0,0);
		(Amult[17] => Cmult[56]) = (0,0);
		(Amult[18] => Cmult[56]) = (0,0);
		(Amult[19] => Cmult[56]) = (0,0);
		(Amult[20] => Cmult[56]) = (0,0);
		(Amult[21] => Cmult[56]) = (0,0);
		(Amult[22] => Cmult[56]) = (0,0);
		(Amult[23] => Cmult[56]) = (0,0);
		(Amult[24] => Cmult[56]) = (0,0);
		(Amult[25] => Cmult[56]) = (0,0);
		(Amult[26] => Cmult[56]) = (0,0);
		(Amult[27] => Cmult[56]) = (0,0);
		(Amult[28] => Cmult[56]) = (0,0);
		(Amult[29] => Cmult[56]) = (0,0);
		(Amult[30] => Cmult[56]) = (0,0);
		(Amult[31] => Cmult[56]) = (0,0);
		(Bmult[0]  => Cmult[56]) = (0,0);
		(Bmult[1]  => Cmult[56]) = (0,0);
		(Bmult[2]  => Cmult[56]) = (0,0);
		(Bmult[3]  => Cmult[56]) = (0,0);
		(Bmult[4]  => Cmult[56]) = (0,0);
		(Bmult[5]  => Cmult[56]) = (0,0);
		(Bmult[6]  => Cmult[56]) = (0,0);
		(Bmult[7]  => Cmult[56]) = (0,0);
		(Bmult[8]  => Cmult[56]) = (0,0);
		(Bmult[9]  => Cmult[56]) = (0,0);
		(Bmult[10] => Cmult[56]) = (0,0);
		(Bmult[11] => Cmult[56]) = (0,0);
		(Bmult[12] => Cmult[56]) = (0,0);
		(Bmult[13] => Cmult[56]) = (0,0);
		(Bmult[14] => Cmult[56]) = (0,0);
		(Bmult[15] => Cmult[56]) = (0,0);
		(Bmult[16] => Cmult[56]) = (0,0);
		(Bmult[17] => Cmult[56]) = (0,0);
		(Bmult[18] => Cmult[56]) = (0,0);
		(Bmult[19] => Cmult[56]) = (0,0);
		(Bmult[20] => Cmult[56]) = (0,0);
		(Bmult[21] => Cmult[56]) = (0,0);
		(Bmult[22] => Cmult[56]) = (0,0);
		(Bmult[23] => Cmult[56]) = (0,0);
		(Bmult[24] => Cmult[56]) = (0,0);
		(Bmult[25] => Cmult[56]) = (0,0);
		(Bmult[26] => Cmult[56]) = (0,0);
		(Bmult[27] => Cmult[56]) = (0,0);
		(Bmult[28] => Cmult[56]) = (0,0);
		(Bmult[29] => Cmult[56]) = (0,0);
		(Bmult[30] => Cmult[56]) = (0,0);
		(Bmult[31] => Cmult[56]) = (0,0);		
		(Valid_mult[0] => Cmult[56]) = (0,0);
		(Valid_mult[1] => Cmult[56]) = (0,0);
		(sel_mul_32x32 => Cmult[56]) = (0,0);
		(Amult[0]  => Cmult[57]) = (0,0);
		(Amult[1]  => Cmult[57]) = (0,0);
		(Amult[2]  => Cmult[57]) = (0,0);
		(Amult[3]  => Cmult[57]) = (0,0);
		(Amult[4]  => Cmult[57]) = (0,0);
		(Amult[5]  => Cmult[57]) = (0,0);
		(Amult[6]  => Cmult[57]) = (0,0);
		(Amult[7]  => Cmult[57]) = (0,0);
		(Amult[8]  => Cmult[57]) = (0,0);
		(Amult[9]  => Cmult[57]) = (0,0);
		(Amult[10] => Cmult[57]) = (0,0);
		(Amult[11] => Cmult[57]) = (0,0);
		(Amult[12] => Cmult[57]) = (0,0);
		(Amult[13] => Cmult[57]) = (0,0);
		(Amult[14] => Cmult[57]) = (0,0);
		(Amult[15] => Cmult[57]) = (0,0);
		(Amult[16] => Cmult[57]) = (0,0);
		(Amult[17] => Cmult[57]) = (0,0);
		(Amult[18] => Cmult[57]) = (0,0);
		(Amult[19] => Cmult[57]) = (0,0);
		(Amult[20] => Cmult[57]) = (0,0);
		(Amult[21] => Cmult[57]) = (0,0);
		(Amult[22] => Cmult[57]) = (0,0);
		(Amult[23] => Cmult[57]) = (0,0);
		(Amult[24] => Cmult[57]) = (0,0);
		(Amult[25] => Cmult[57]) = (0,0);
		(Amult[26] => Cmult[57]) = (0,0);
		(Amult[27] => Cmult[57]) = (0,0);
		(Amult[28] => Cmult[57]) = (0,0);
		(Amult[29] => Cmult[57]) = (0,0);
		(Amult[30] => Cmult[57]) = (0,0);
		(Amult[31] => Cmult[57]) = (0,0);
		(Bmult[0]  => Cmult[57]) = (0,0);
		(Bmult[1]  => Cmult[57]) = (0,0);
		(Bmult[2]  => Cmult[57]) = (0,0);
		(Bmult[3]  => Cmult[57]) = (0,0);
		(Bmult[4]  => Cmult[57]) = (0,0);
		(Bmult[5]  => Cmult[57]) = (0,0);
		(Bmult[6]  => Cmult[57]) = (0,0);
		(Bmult[7]  => Cmult[57]) = (0,0);
		(Bmult[8]  => Cmult[57]) = (0,0);
		(Bmult[9]  => Cmult[57]) = (0,0);
		(Bmult[10] => Cmult[57]) = (0,0);
		(Bmult[11] => Cmult[57]) = (0,0);
		(Bmult[12] => Cmult[57]) = (0,0);
		(Bmult[13] => Cmult[57]) = (0,0);
		(Bmult[14] => Cmult[57]) = (0,0);
		(Bmult[15] => Cmult[57]) = (0,0);
		(Bmult[16] => Cmult[57]) = (0,0);
		(Bmult[17] => Cmult[57]) = (0,0);
		(Bmult[18] => Cmult[57]) = (0,0);
		(Bmult[19] => Cmult[57]) = (0,0);
		(Bmult[20] => Cmult[57]) = (0,0);
		(Bmult[21] => Cmult[57]) = (0,0);
		(Bmult[22] => Cmult[57]) = (0,0);
		(Bmult[23] => Cmult[57]) = (0,0);
		(Bmult[24] => Cmult[57]) = (0,0);
		(Bmult[25] => Cmult[57]) = (0,0);
		(Bmult[26] => Cmult[57]) = (0,0);
		(Bmult[27] => Cmult[57]) = (0,0);
		(Bmult[28] => Cmult[57]) = (0,0);
		(Bmult[29] => Cmult[57]) = (0,0);
		(Bmult[30] => Cmult[57]) = (0,0);
		(Bmult[31] => Cmult[57]) = (0,0);		
		(Valid_mult[0] => Cmult[57]) = (0,0);
		(Valid_mult[1] => Cmult[57]) = (0,0);
		(sel_mul_32x32 => Cmult[57]) = (0,0);
		(Amult[0]  => Cmult[58]) = (0,0);
		(Amult[1]  => Cmult[58]) = (0,0);
		(Amult[2]  => Cmult[58]) = (0,0);
		(Amult[3]  => Cmult[58]) = (0,0);
		(Amult[4]  => Cmult[58]) = (0,0);
		(Amult[5]  => Cmult[58]) = (0,0);
		(Amult[6]  => Cmult[58]) = (0,0);
		(Amult[7]  => Cmult[58]) = (0,0);
		(Amult[8]  => Cmult[58]) = (0,0);
		(Amult[9]  => Cmult[58]) = (0,0);
		(Amult[10] => Cmult[58]) = (0,0);
		(Amult[11] => Cmult[58]) = (0,0);
		(Amult[12] => Cmult[58]) = (0,0);
		(Amult[13] => Cmult[58]) = (0,0);
		(Amult[14] => Cmult[58]) = (0,0);
		(Amult[15] => Cmult[58]) = (0,0);
		(Amult[16] => Cmult[58]) = (0,0);
		(Amult[17] => Cmult[58]) = (0,0);
		(Amult[18] => Cmult[58]) = (0,0);
		(Amult[19] => Cmult[58]) = (0,0);
		(Amult[20] => Cmult[58]) = (0,0);
		(Amult[21] => Cmult[58]) = (0,0);
		(Amult[22] => Cmult[58]) = (0,0);
		(Amult[23] => Cmult[58]) = (0,0);
		(Amult[24] => Cmult[58]) = (0,0);
		(Amult[25] => Cmult[58]) = (0,0);
		(Amult[26] => Cmult[58]) = (0,0);
		(Amult[27] => Cmult[58]) = (0,0);
		(Amult[28] => Cmult[58]) = (0,0);
		(Amult[29] => Cmult[58]) = (0,0);
		(Amult[30] => Cmult[58]) = (0,0);
		(Amult[31] => Cmult[58]) = (0,0);
		(Bmult[0]  => Cmult[58]) = (0,0);
		(Bmult[1]  => Cmult[58]) = (0,0);
		(Bmult[2]  => Cmult[58]) = (0,0);
		(Bmult[3]  => Cmult[58]) = (0,0);
		(Bmult[4]  => Cmult[58]) = (0,0);
		(Bmult[5]  => Cmult[58]) = (0,0);
		(Bmult[6]  => Cmult[58]) = (0,0);
		(Bmult[7]  => Cmult[58]) = (0,0);
		(Bmult[8]  => Cmult[58]) = (0,0);
		(Bmult[9]  => Cmult[58]) = (0,0);
		(Bmult[10] => Cmult[58]) = (0,0);
		(Bmult[11] => Cmult[58]) = (0,0);
		(Bmult[12] => Cmult[58]) = (0,0);
		(Bmult[13] => Cmult[58]) = (0,0);
		(Bmult[14] => Cmult[58]) = (0,0);
		(Bmult[15] => Cmult[58]) = (0,0);
		(Bmult[16] => Cmult[58]) = (0,0);
		(Bmult[17] => Cmult[58]) = (0,0);
		(Bmult[18] => Cmult[58]) = (0,0);
		(Bmult[19] => Cmult[58]) = (0,0);
		(Bmult[20] => Cmult[58]) = (0,0);
		(Bmult[21] => Cmult[58]) = (0,0);
		(Bmult[22] => Cmult[58]) = (0,0);
		(Bmult[23] => Cmult[58]) = (0,0);
		(Bmult[24] => Cmult[58]) = (0,0);
		(Bmult[25] => Cmult[58]) = (0,0);
		(Bmult[26] => Cmult[58]) = (0,0);
		(Bmult[27] => Cmult[58]) = (0,0);
		(Bmult[28] => Cmult[58]) = (0,0);
		(Bmult[29] => Cmult[58]) = (0,0);
		(Bmult[30] => Cmult[58]) = (0,0);
		(Bmult[31] => Cmult[58]) = (0,0);		
		(Valid_mult[0] => Cmult[58]) = (0,0);
		(Valid_mult[1] => Cmult[58]) = (0,0);
		(sel_mul_32x32 => Cmult[58]) = (0,0);	
		(Amult[0]  => Cmult[59]) = (0,0);
		(Amult[1]  => Cmult[59]) = (0,0);
		(Amult[2]  => Cmult[59]) = (0,0);
		(Amult[3]  => Cmult[59]) = (0,0);
		(Amult[4]  => Cmult[59]) = (0,0);
		(Amult[5]  => Cmult[59]) = (0,0);
		(Amult[6]  => Cmult[59]) = (0,0);
		(Amult[7]  => Cmult[59]) = (0,0);
		(Amult[8]  => Cmult[59]) = (0,0);
		(Amult[9]  => Cmult[59]) = (0,0);
		(Amult[10] => Cmult[59]) = (0,0);
		(Amult[11] => Cmult[59]) = (0,0);
		(Amult[12] => Cmult[59]) = (0,0);
		(Amult[13] => Cmult[59]) = (0,0);
		(Amult[14] => Cmult[59]) = (0,0);
		(Amult[15] => Cmult[59]) = (0,0);
		(Amult[16] => Cmult[59]) = (0,0);
		(Amult[17] => Cmult[59]) = (0,0);
		(Amult[18] => Cmult[59]) = (0,0);
		(Amult[19] => Cmult[59]) = (0,0);
		(Amult[20] => Cmult[59]) = (0,0);
		(Amult[21] => Cmult[59]) = (0,0);
		(Amult[22] => Cmult[59]) = (0,0);
		(Amult[23] => Cmult[59]) = (0,0);
		(Amult[24] => Cmult[59]) = (0,0);
		(Amult[25] => Cmult[59]) = (0,0);
		(Amult[26] => Cmult[59]) = (0,0);
		(Amult[27] => Cmult[59]) = (0,0);
		(Amult[28] => Cmult[59]) = (0,0);
		(Amult[29] => Cmult[59]) = (0,0);
		(Amult[30] => Cmult[59]) = (0,0);
		(Amult[31] => Cmult[59]) = (0,0);
		(Bmult[0]  => Cmult[59]) = (0,0);
		(Bmult[1]  => Cmult[59]) = (0,0);
		(Bmult[2]  => Cmult[59]) = (0,0);
		(Bmult[3]  => Cmult[59]) = (0,0);
		(Bmult[4]  => Cmult[59]) = (0,0);
		(Bmult[5]  => Cmult[59]) = (0,0);
		(Bmult[6]  => Cmult[59]) = (0,0);
		(Bmult[7]  => Cmult[59]) = (0,0);
		(Bmult[8]  => Cmult[59]) = (0,0);
		(Bmult[9]  => Cmult[59]) = (0,0);
		(Bmult[10] => Cmult[59]) = (0,0);
		(Bmult[11] => Cmult[59]) = (0,0);
		(Bmult[12] => Cmult[59]) = (0,0);
		(Bmult[13] => Cmult[59]) = (0,0);
		(Bmult[14] => Cmult[59]) = (0,0);
		(Bmult[15] => Cmult[59]) = (0,0);
		(Bmult[16] => Cmult[59]) = (0,0);
		(Bmult[17] => Cmult[59]) = (0,0);
		(Bmult[18] => Cmult[59]) = (0,0);
		(Bmult[19] => Cmult[59]) = (0,0);
		(Bmult[20] => Cmult[59]) = (0,0);
		(Bmult[21] => Cmult[59]) = (0,0);
		(Bmult[22] => Cmult[59]) = (0,0);
		(Bmult[23] => Cmult[59]) = (0,0);
		(Bmult[24] => Cmult[59]) = (0,0);
		(Bmult[25] => Cmult[59]) = (0,0);
		(Bmult[26] => Cmult[59]) = (0,0);
		(Bmult[27] => Cmult[59]) = (0,0);
		(Bmult[28] => Cmult[59]) = (0,0);
		(Bmult[29] => Cmult[59]) = (0,0);
		(Bmult[30] => Cmult[59]) = (0,0);
		(Bmult[31] => Cmult[59]) = (0,0);		
		(Valid_mult[0] => Cmult[59]) = (0,0);
		(Valid_mult[1] => Cmult[59]) = (0,0);
		(sel_mul_32x32 => Cmult[59]) = (0,0);
		(Amult[0]  => Cmult[60]) = (0,0);
		(Amult[1]  => Cmult[60]) = (0,0);
		(Amult[2]  => Cmult[60]) = (0,0);
		(Amult[3]  => Cmult[60]) = (0,0);
		(Amult[4]  => Cmult[60]) = (0,0);
		(Amult[5]  => Cmult[60]) = (0,0);
		(Amult[6]  => Cmult[60]) = (0,0);
		(Amult[7]  => Cmult[60]) = (0,0);
		(Amult[8]  => Cmult[60]) = (0,0);
		(Amult[9]  => Cmult[60]) = (0,0);
		(Amult[10] => Cmult[60]) = (0,0);
		(Amult[11] => Cmult[60]) = (0,0);
		(Amult[12] => Cmult[60]) = (0,0);
		(Amult[13] => Cmult[60]) = (0,0);
		(Amult[14] => Cmult[60]) = (0,0);
		(Amult[15] => Cmult[60]) = (0,0);
		(Amult[16] => Cmult[60]) = (0,0);
		(Amult[17] => Cmult[60]) = (0,0);
		(Amult[18] => Cmult[60]) = (0,0);
		(Amult[19] => Cmult[60]) = (0,0);
		(Amult[20] => Cmult[60]) = (0,0);
		(Amult[21] => Cmult[60]) = (0,0);
		(Amult[22] => Cmult[60]) = (0,0);
		(Amult[23] => Cmult[60]) = (0,0);
		(Amult[24] => Cmult[60]) = (0,0);
		(Amult[25] => Cmult[60]) = (0,0);
		(Amult[26] => Cmult[60]) = (0,0);
		(Amult[27] => Cmult[60]) = (0,0);
		(Amult[28] => Cmult[60]) = (0,0);
		(Amult[29] => Cmult[60]) = (0,0);
		(Amult[30] => Cmult[60]) = (0,0);
		(Amult[31] => Cmult[60]) = (0,0);
		(Bmult[0]  => Cmult[60]) = (0,0);
		(Bmult[1]  => Cmult[60]) = (0,0);
		(Bmult[2]  => Cmult[60]) = (0,0);
		(Bmult[3]  => Cmult[60]) = (0,0);
		(Bmult[4]  => Cmult[60]) = (0,0);
		(Bmult[5]  => Cmult[60]) = (0,0);
		(Bmult[6]  => Cmult[60]) = (0,0);
		(Bmult[7]  => Cmult[60]) = (0,0);
		(Bmult[8]  => Cmult[60]) = (0,0);
		(Bmult[9]  => Cmult[60]) = (0,0);
		(Bmult[10] => Cmult[60]) = (0,0);
		(Bmult[11] => Cmult[60]) = (0,0);
		(Bmult[12] => Cmult[60]) = (0,0);
		(Bmult[13] => Cmult[60]) = (0,0);
		(Bmult[14] => Cmult[60]) = (0,0);
		(Bmult[15] => Cmult[60]) = (0,0);
		(Bmult[16] => Cmult[60]) = (0,0);
		(Bmult[17] => Cmult[60]) = (0,0);
		(Bmult[18] => Cmult[60]) = (0,0);
		(Bmult[19] => Cmult[60]) = (0,0);
		(Bmult[20] => Cmult[60]) = (0,0);
		(Bmult[21] => Cmult[60]) = (0,0);
		(Bmult[22] => Cmult[60]) = (0,0);
		(Bmult[23] => Cmult[60]) = (0,0);
		(Bmult[24] => Cmult[60]) = (0,0);
		(Bmult[25] => Cmult[60]) = (0,0);
		(Bmult[26] => Cmult[60]) = (0,0);
		(Bmult[27] => Cmult[60]) = (0,0);
		(Bmult[28] => Cmult[60]) = (0,0);
		(Bmult[29] => Cmult[60]) = (0,0);
		(Bmult[30] => Cmult[60]) = (0,0);
		(Bmult[31] => Cmult[60]) = (0,0);		
		(Valid_mult[0] => Cmult[60]) = (0,0);
		(Valid_mult[1] => Cmult[60]) = (0,0);
		(sel_mul_32x32 => Cmult[60]) = (0,0);
		(Amult[0]  => Cmult[61]) = (0,0);
		(Amult[1]  => Cmult[61]) = (0,0);
		(Amult[2]  => Cmult[61]) = (0,0);
		(Amult[3]  => Cmult[61]) = (0,0);
		(Amult[4]  => Cmult[61]) = (0,0);
		(Amult[5]  => Cmult[61]) = (0,0);
		(Amult[6]  => Cmult[61]) = (0,0);
		(Amult[7]  => Cmult[61]) = (0,0);
		(Amult[8]  => Cmult[61]) = (0,0);
		(Amult[9]  => Cmult[61]) = (0,0);
		(Amult[10] => Cmult[61]) = (0,0);
		(Amult[11] => Cmult[61]) = (0,0);
		(Amult[12] => Cmult[61]) = (0,0);
		(Amult[13] => Cmult[61]) = (0,0);
		(Amult[14] => Cmult[61]) = (0,0);
		(Amult[15] => Cmult[61]) = (0,0);
		(Amult[16] => Cmult[61]) = (0,0);
		(Amult[17] => Cmult[61]) = (0,0);
		(Amult[18] => Cmult[61]) = (0,0);
		(Amult[19] => Cmult[61]) = (0,0);
		(Amult[20] => Cmult[61]) = (0,0);
		(Amult[21] => Cmult[61]) = (0,0);
		(Amult[22] => Cmult[61]) = (0,0);
		(Amult[23] => Cmult[61]) = (0,0);
		(Amult[24] => Cmult[61]) = (0,0);
		(Amult[25] => Cmult[61]) = (0,0);
		(Amult[26] => Cmult[61]) = (0,0);
		(Amult[27] => Cmult[61]) = (0,0);
		(Amult[28] => Cmult[61]) = (0,0);
		(Amult[29] => Cmult[61]) = (0,0);
		(Amult[30] => Cmult[61]) = (0,0);
		(Amult[31] => Cmult[61]) = (0,0);
		(Bmult[0]  => Cmult[61]) = (0,0);
		(Bmult[1]  => Cmult[61]) = (0,0);
		(Bmult[2]  => Cmult[61]) = (0,0);
		(Bmult[3]  => Cmult[61]) = (0,0);
		(Bmult[4]  => Cmult[61]) = (0,0);
		(Bmult[5]  => Cmult[61]) = (0,0);
		(Bmult[6]  => Cmult[61]) = (0,0);
		(Bmult[7]  => Cmult[61]) = (0,0);
		(Bmult[8]  => Cmult[61]) = (0,0);
		(Bmult[9]  => Cmult[61]) = (0,0);
		(Bmult[10] => Cmult[61]) = (0,0);
		(Bmult[11] => Cmult[61]) = (0,0);
		(Bmult[12] => Cmult[61]) = (0,0);
		(Bmult[13] => Cmult[61]) = (0,0);
		(Bmult[14] => Cmult[61]) = (0,0);
		(Bmult[15] => Cmult[61]) = (0,0);
		(Bmult[16] => Cmult[61]) = (0,0);
		(Bmult[17] => Cmult[61]) = (0,0);
		(Bmult[18] => Cmult[61]) = (0,0);
		(Bmult[19] => Cmult[61]) = (0,0);
		(Bmult[20] => Cmult[61]) = (0,0);
		(Bmult[21] => Cmult[61]) = (0,0);
		(Bmult[22] => Cmult[61]) = (0,0);
		(Bmult[23] => Cmult[61]) = (0,0);
		(Bmult[24] => Cmult[61]) = (0,0);
		(Bmult[25] => Cmult[61]) = (0,0);
		(Bmult[26] => Cmult[61]) = (0,0);
		(Bmult[27] => Cmult[61]) = (0,0);
		(Bmult[28] => Cmult[61]) = (0,0);
		(Bmult[29] => Cmult[61]) = (0,0);
		(Bmult[30] => Cmult[61]) = (0,0);
		(Bmult[31] => Cmult[61]) = (0,0);		
		(Valid_mult[0] => Cmult[61]) = (0,0);
		(Valid_mult[1] => Cmult[61]) = (0,0);
		(sel_mul_32x32 => Cmult[61]) = (0,0);
		(Amult[0]  => Cmult[62]) = (0,0);
		(Amult[1]  => Cmult[62]) = (0,0);
		(Amult[2]  => Cmult[62]) = (0,0);
		(Amult[3]  => Cmult[62]) = (0,0);
		(Amult[4]  => Cmult[62]) = (0,0);
		(Amult[5]  => Cmult[62]) = (0,0);
		(Amult[6]  => Cmult[62]) = (0,0);
		(Amult[7]  => Cmult[62]) = (0,0);
		(Amult[8]  => Cmult[62]) = (0,0);
		(Amult[9]  => Cmult[62]) = (0,0);
		(Amult[10] => Cmult[62]) = (0,0);
		(Amult[11] => Cmult[62]) = (0,0);
		(Amult[12] => Cmult[62]) = (0,0);
		(Amult[13] => Cmult[62]) = (0,0);
		(Amult[14] => Cmult[62]) = (0,0);
		(Amult[15] => Cmult[62]) = (0,0);
		(Amult[16] => Cmult[62]) = (0,0);
		(Amult[17] => Cmult[62]) = (0,0);
		(Amult[18] => Cmult[62]) = (0,0);
		(Amult[19] => Cmult[62]) = (0,0);
		(Amult[20] => Cmult[62]) = (0,0);
		(Amult[21] => Cmult[62]) = (0,0);
		(Amult[22] => Cmult[62]) = (0,0);
		(Amult[23] => Cmult[62]) = (0,0);
		(Amult[24] => Cmult[62]) = (0,0);
		(Amult[25] => Cmult[62]) = (0,0);
		(Amult[26] => Cmult[62]) = (0,0);
		(Amult[27] => Cmult[62]) = (0,0);
		(Amult[28] => Cmult[62]) = (0,0);
		(Amult[29] => Cmult[62]) = (0,0);
		(Amult[30] => Cmult[62]) = (0,0);
		(Amult[31] => Cmult[62]) = (0,0);
		(Bmult[0]  => Cmult[62]) = (0,0);
		(Bmult[1]  => Cmult[62]) = (0,0);
		(Bmult[2]  => Cmult[62]) = (0,0);
		(Bmult[3]  => Cmult[62]) = (0,0);
		(Bmult[4]  => Cmult[62]) = (0,0);
		(Bmult[5]  => Cmult[62]) = (0,0);
		(Bmult[6]  => Cmult[62]) = (0,0);
		(Bmult[7]  => Cmult[62]) = (0,0);
		(Bmult[8]  => Cmult[62]) = (0,0);
		(Bmult[9]  => Cmult[62]) = (0,0);
		(Bmult[10] => Cmult[62]) = (0,0);
		(Bmult[11] => Cmult[62]) = (0,0);
		(Bmult[12] => Cmult[62]) = (0,0);
		(Bmult[13] => Cmult[62]) = (0,0);
		(Bmult[14] => Cmult[62]) = (0,0);
		(Bmult[15] => Cmult[62]) = (0,0);
		(Bmult[16] => Cmult[62]) = (0,0);
		(Bmult[17] => Cmult[62]) = (0,0);
		(Bmult[18] => Cmult[62]) = (0,0);
		(Bmult[19] => Cmult[62]) = (0,0);
		(Bmult[20] => Cmult[62]) = (0,0);
		(Bmult[21] => Cmult[62]) = (0,0);
		(Bmult[22] => Cmult[62]) = (0,0);
		(Bmult[23] => Cmult[62]) = (0,0);
		(Bmult[24] => Cmult[62]) = (0,0);
		(Bmult[25] => Cmult[62]) = (0,0);
		(Bmult[26] => Cmult[62]) = (0,0);
		(Bmult[27] => Cmult[62]) = (0,0);
		(Bmult[28] => Cmult[62]) = (0,0);
		(Bmult[29] => Cmult[62]) = (0,0);
		(Bmult[30] => Cmult[62]) = (0,0);
		(Bmult[31] => Cmult[62]) = (0,0);		
		(Valid_mult[0] => Cmult[62]) = (0,0);
		(Valid_mult[1] => Cmult[62]) = (0,0);
		(sel_mul_32x32 => Cmult[62]) = (0,0);
		(Amult[0]  => Cmult[63]) = (0,0);
		(Amult[1]  => Cmult[63]) = (0,0);
		(Amult[2]  => Cmult[63]) = (0,0);
		(Amult[3]  => Cmult[63]) = (0,0);
		(Amult[4]  => Cmult[63]) = (0,0);
		(Amult[5]  => Cmult[63]) = (0,0);
		(Amult[6]  => Cmult[63]) = (0,0);
		(Amult[7]  => Cmult[63]) = (0,0);
		(Amult[8]  => Cmult[63]) = (0,0);
		(Amult[9]  => Cmult[63]) = (0,0);
		(Amult[10] => Cmult[63]) = (0,0);
		(Amult[11] => Cmult[63]) = (0,0);
		(Amult[12] => Cmult[63]) = (0,0);
		(Amult[13] => Cmult[63]) = (0,0);
		(Amult[14] => Cmult[63]) = (0,0);
		(Amult[15] => Cmult[63]) = (0,0);
		(Amult[16] => Cmult[63]) = (0,0);
		(Amult[17] => Cmult[63]) = (0,0);
		(Amult[18] => Cmult[63]) = (0,0);
		(Amult[19] => Cmult[63]) = (0,0);
		(Amult[20] => Cmult[63]) = (0,0);
		(Amult[21] => Cmult[63]) = (0,0);
		(Amult[22] => Cmult[63]) = (0,0);
		(Amult[23] => Cmult[63]) = (0,0);
		(Amult[24] => Cmult[63]) = (0,0);
		(Amult[25] => Cmult[63]) = (0,0);
		(Amult[26] => Cmult[63]) = (0,0);
		(Amult[27] => Cmult[63]) = (0,0);
		(Amult[28] => Cmult[63]) = (0,0);
		(Amult[29] => Cmult[63]) = (0,0);
		(Amult[30] => Cmult[63]) = (0,0);
		(Amult[31] => Cmult[63]) = (0,0);
		(Bmult[0]  => Cmult[63]) = (0,0);
		(Bmult[1]  => Cmult[63]) = (0,0);
		(Bmult[2]  => Cmult[63]) = (0,0);
		(Bmult[3]  => Cmult[63]) = (0,0);
		(Bmult[4]  => Cmult[63]) = (0,0);
		(Bmult[5]  => Cmult[63]) = (0,0);
		(Bmult[6]  => Cmult[63]) = (0,0);
		(Bmult[7]  => Cmult[63]) = (0,0);
		(Bmult[8]  => Cmult[63]) = (0,0);
		(Bmult[9]  => Cmult[63]) = (0,0);
		(Bmult[10] => Cmult[63]) = (0,0);
		(Bmult[11] => Cmult[63]) = (0,0);
		(Bmult[12] => Cmult[63]) = (0,0);
		(Bmult[13] => Cmult[63]) = (0,0);
		(Bmult[14] => Cmult[63]) = (0,0);
		(Bmult[15] => Cmult[63]) = (0,0);
		(Bmult[16] => Cmult[63]) = (0,0);
		(Bmult[17] => Cmult[63]) = (0,0);
		(Bmult[18] => Cmult[63]) = (0,0);
		(Bmult[19] => Cmult[63]) = (0,0);
		(Bmult[20] => Cmult[63]) = (0,0);
		(Bmult[21] => Cmult[63]) = (0,0);
		(Bmult[22] => Cmult[63]) = (0,0);
		(Bmult[23] => Cmult[63]) = (0,0);
		(Bmult[24] => Cmult[63]) = (0,0);
		(Bmult[25] => Cmult[63]) = (0,0);
		(Bmult[26] => Cmult[63]) = (0,0);
		(Bmult[27] => Cmult[63]) = (0,0);
		(Bmult[28] => Cmult[63]) = (0,0);
		(Bmult[29] => Cmult[63]) = (0,0);
		(Bmult[30] => Cmult[63]) = (0,0);
		(Bmult[31] => Cmult[63]) = (0,0);		
		(Valid_mult[0] => Cmult[63]) = (0,0);
		(Valid_mult[1] => Cmult[63]) = (0,0);
		(sel_mul_32x32 => Cmult[63]) = (0,0);		
    endspecify
`endif
	
	always @(*) begin
		if (sel_mul_32x32 == 1'b1) begin
			if (Valid_mult[0] == 1'b1) begin
				Cmult <= Amult * Bmult;
			end
		end else begin
			if (Valid_mult[0] == 1'b1) begin
				Cmult[31:0] <= Amult[15:0] * Bmult[15:0];
			end
			if (Valid_mult[1] == 1'b1) begin
				Cmult[63:32] <= Amult[31:16] * Bmult[31:16];
			end
		end
	end


endmodule
// ../../../quicklogic/pp3/primitives/mult/mult.sim.v }}}

// ../../../quicklogic/pp3/primitives/gmux/gmux_ip.sim.v {{{
(* whitebox *)
module GMUX_IP (IP, IC, IS0, IZ);

    input  wire IP;
    input  wire IC;
    input  wire IS0;

    (* clkbuf_driver *)
    output wire IZ;

    specify
        (IP => IZ) = (0,0);
		(IC => IZ) = (0,0);
		(IS0 => IZ) = (0,0);
    endspecify

    assign IZ = IS0 ? IC : IP;

endmodule
// ../../../quicklogic/pp3/primitives/gmux/gmux_ip.sim.v }}}

// ../../../quicklogic/pp3/primitives/gmux/gmux_ic.sim.v {{{
(* whitebox *)
module GMUX_IC (IC, IS0, IZ);

    input  wire IC;
    input  wire IS0;

    (* clkbuf_driver *)
    output wire IZ;
	
    specify
        (IC => IZ) = (0,0);
		(IS0 => IZ) = (0,0);
    endspecify

    assign IZ = IS0 ? IC : 1'bx;

endmodule
// ../../../quicklogic/pp3/primitives/gmux/gmux_ic.sim.v }}}
