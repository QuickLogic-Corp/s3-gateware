//`include "C:/QuickLogic/QuickWorks_2016.2_Release/spde/data/PolarPro-III/AL4S3B/rrw/fifo_blk.v" 
`ifdef f512x8_512x8
`else
`define f512x8_512x8
/************************************************************************
** File : f512x8_512x8.v
** Design Date: July 18,2012
** Creation Date: Wed May 13 16:02:49 2020

** Created By SpDE Version: SpDE 2016.2 Release
** Author: QuickLogic Corporation,
** Copyright (C) 1998, Customers of QuickLogic may copy and modify this
** file for use in designing QuickLogic devices only.
** Description : This file is autogenerated RTL code that describes the
** top level design for FIFO using QuickLogic's
** RAM block resources.
************************************************************************/
module f512x8_512x8(DIN,Fifo_Push_Flush,Fifo_Pop_Flush,PUSH,POP,Clk,
       Clk_En,Fifo_Dir,Async_Flush,
       Almost_Full,Almost_Empty,PUSH_FLAG,POP_FLAG,DOUT);


input Fifo_Push_Flush,Fifo_Pop_Flush;
input Clk;
input PUSH,POP;
input [7:0] DIN;
input Clk_En,Fifo_Dir,Async_Flush;
output [7:0] DOUT;
output [3:0] PUSH_FLAG,POP_FLAG;
output Almost_Full,Almost_Empty;

parameter wr_depth_int = 512;
parameter rd_depth_int = 512;
parameter wr_width_int = 8;
parameter rd_width_int = 8;
parameter reg_rd_int = 0;
parameter sync_fifo_int = 1;

parameter data_depth_int = 512;
parameter data_width_int = 8;

supply0 GND;
supply1 VCC;
//FIFO
FIFO_8K_BLK
#(
//    wr_depth_int, rd_depth_int,
//    wr_width_int,rd_width_int,
    .data_depth_int(data_depth_int),
    .data_width_int(data_width_int),
    .reg_rd_int(reg_rd_int),
    .sync_fifo_int(sync_fifo_int)) 
FIFO_INST (.DIN(DIN),.PUSH(PUSH),.POP(POP),.Fifo_Push_Flush(Fifo_Push_Flush),.Fifo_Pop_Flush(Fifo_Pop_Flush),
           .Push_Clk(Clk),.Pop_Clk(Clk),.PUSH_FLAG(PUSH_FLAG),.POP_FLAG(POP_FLAG),
      .Push_Clk_En(Clk_En),.Pop_Clk_En(Clk_En),.Fifo_Dir(Fifo_Dir),.Async_Flush(Async_Flush),
//      .Push_Clk_Sel(GND),
//      .Pop_Clk_Sel(GND),
//      .Async_Flush_Sel(GND),
           .Almost_Full(Almost_Full),.Almost_Empty(Almost_Empty),.DOUT(DOUT)
//           ,
//        .LS(1'b0), .SD(1'b0), .DS(1'b0), .LS_RB1(1'b0), .SD_RB1(1'b0), .DS_RB1(1'b0)
    );
endmodule
`endif
